library ieee;
use ieee.std_logic_1164.all;

package liaison_tb_data is

    constant count : integer := 256;

    type inputvect_t is array(0 to count-1, 0 to 4) of std_logic_vector(7 downto 0);
    type outputvect_t is array(0 to count-1) of std_logic_vector(14 downto 0);

    -- 0 => (0 => "00000000", 1 => "00000000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
    constant input : inputvect_t := (
            0 => (0 => "00000000", 1 => "00000000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            1 => (0 => "00000001", 1 => "00000001", 2 => "00000001", 3 => "00000001", 4 => "00000000"),
            2 => (0 => "00000010", 1 => "00000010", 2 => "00000010", 3 => "00000010", 4 => "00000000"),
            3 => (0 => "00000011", 1 => "00000011", 2 => "00000011", 3 => "00000011", 4 => "00000000"),
            4 => (0 => "00000100", 1 => "00000100", 2 => "00000100", 3 => "00000100", 4 => "00000000"),
            5 => (0 => "00000101", 1 => "00000101", 2 => "00000101", 3 => "00000101", 4 => "00000000"),
            6 => (0 => "00000110", 1 => "00000110", 2 => "00000110", 3 => "00000110", 4 => "00000000"),
            7 => (0 => "00000111", 1 => "00000111", 2 => "00000111", 3 => "00000111", 4 => "00000000"),
            8 => (0 => "00001000", 1 => "00001000", 2 => "00001000", 3 => "00001000", 4 => "00000000"),
            9 => (0 => "00001001", 1 => "00001001", 2 => "00001001", 3 => "00001001", 4 => "00000000"),
            10 => (0 => "00001010", 1 => "00001010", 2 => "00001010", 3 => "00001010", 4 => "00000000"),
            11 => (0 => "00001011", 1 => "00001011", 2 => "00001011", 3 => "00001011", 4 => "00000000"),
            12 => (0 => "00001100", 1 => "00001100", 2 => "00001100", 3 => "00001100", 4 => "00000000"),
            13 => (0 => "00001101", 1 => "00001101", 2 => "00001101", 3 => "00001101", 4 => "00000000"),
            14 => (0 => "00001110", 1 => "00001110", 2 => "00001110", 3 => "00001110", 4 => "00000000"),
            15 => (0 => "00001111", 1 => "00001111", 2 => "00001111", 3 => "00001111", 4 => "00000000"),
            16 => (0 => "00010000", 1 => "00010000", 2 => "00010000", 3 => "00010000", 4 => "00000000"),
            17 => (0 => "00010001", 1 => "00010001", 2 => "00010001", 3 => "00010001", 4 => "00000000"),
            18 => (0 => "00010010", 1 => "00010010", 2 => "00010010", 3 => "00010010", 4 => "00000000"),
            19 => (0 => "00010011", 1 => "00010011", 2 => "00010011", 3 => "00010011", 4 => "00000000"),
            20 => (0 => "00010100", 1 => "00010100", 2 => "00010100", 3 => "00010100", 4 => "00000000"),
            21 => (0 => "00010101", 1 => "00010101", 2 => "00010101", 3 => "00010101", 4 => "00000000"),
            22 => (0 => "00010110", 1 => "00010110", 2 => "00010110", 3 => "00010110", 4 => "00000000"),
            23 => (0 => "00010111", 1 => "00010111", 2 => "00010111", 3 => "00010111", 4 => "00000000"),
            24 => (0 => "00011000", 1 => "00011000", 2 => "00011000", 3 => "00011000", 4 => "00000000"),
            25 => (0 => "00011001", 1 => "00011001", 2 => "00011001", 3 => "00011001", 4 => "00000000"),
            26 => (0 => "00011010", 1 => "00011010", 2 => "00011010", 3 => "00011010", 4 => "00000000"),
            27 => (0 => "00011011", 1 => "00011011", 2 => "00011011", 3 => "00011011", 4 => "00000000"),
            28 => (0 => "00011100", 1 => "00011100", 2 => "00011100", 3 => "00011100", 4 => "00000000"),
            29 => (0 => "00011101", 1 => "00011101", 2 => "00011101", 3 => "00011101", 4 => "00000000"),
            30 => (0 => "00011110", 1 => "00011110", 2 => "00011110", 3 => "00011110", 4 => "00000000"),
            31 => (0 => "00011111", 1 => "00011111", 2 => "00011111", 3 => "00011111", 4 => "00000000"),
            32 => (0 => "00100000", 1 => "00100000", 2 => "00100000", 3 => "00100000", 4 => "00000000"),
            33 => (0 => "00100001", 1 => "00100001", 2 => "00100001", 3 => "00100001", 4 => "00000000"),
            34 => (0 => "00100010", 1 => "00100010", 2 => "00100010", 3 => "00100010", 4 => "00000000"),
            35 => (0 => "00100011", 1 => "00100011", 2 => "00100011", 3 => "00100011", 4 => "00000000"),
            36 => (0 => "00100100", 1 => "00100100", 2 => "00100100", 3 => "00100100", 4 => "00000000"),
            37 => (0 => "00100101", 1 => "00100101", 2 => "00100101", 3 => "00100101", 4 => "00000000"),
            38 => (0 => "00100110", 1 => "00100110", 2 => "00100110", 3 => "00100110", 4 => "00000000"),
            39 => (0 => "00100111", 1 => "00100111", 2 => "00100111", 3 => "00100111", 4 => "00000000"),
            40 => (0 => "00101000", 1 => "00101000", 2 => "00101000", 3 => "00101000", 4 => "00000000"),
            41 => (0 => "00101001", 1 => "00101001", 2 => "00101001", 3 => "00101001", 4 => "00000000"),
            42 => (0 => "00101010", 1 => "00101010", 2 => "00101010", 3 => "00101010", 4 => "00000000"),
            43 => (0 => "00101011", 1 => "00101011", 2 => "00101011", 3 => "00101011", 4 => "00000000"),
            44 => (0 => "00101100", 1 => "00101100", 2 => "00101100", 3 => "00101100", 4 => "00000000"),
            45 => (0 => "00101101", 1 => "00101101", 2 => "00101101", 3 => "00101101", 4 => "00000000"),
            46 => (0 => "00101110", 1 => "00101110", 2 => "00101110", 3 => "00101110", 4 => "00000000"),
            47 => (0 => "00101111", 1 => "00101111", 2 => "00101111", 3 => "00101111", 4 => "00000000"),
            48 => (0 => "00110000", 1 => "00110000", 2 => "00110000", 3 => "00110000", 4 => "00000000"),
            49 => (0 => "00110001", 1 => "00110001", 2 => "00110001", 3 => "00110001", 4 => "00000000"),
            50 => (0 => "00110010", 1 => "00110010", 2 => "00110010", 3 => "00110010", 4 => "00000000"),
            51 => (0 => "00110011", 1 => "00110011", 2 => "00110011", 3 => "00110011", 4 => "00000000"),
            52 => (0 => "00110100", 1 => "00110100", 2 => "00110100", 3 => "00110100", 4 => "00000000"),
            53 => (0 => "00110101", 1 => "00110101", 2 => "00110101", 3 => "00110101", 4 => "00000000"),
            54 => (0 => "00110110", 1 => "00110110", 2 => "00110110", 3 => "00110110", 4 => "00000000"),
            55 => (0 => "00110111", 1 => "00110111", 2 => "00110111", 3 => "00110111", 4 => "00000000"),
            56 => (0 => "00111000", 1 => "00111000", 2 => "00111000", 3 => "00111000", 4 => "00000000"),
            57 => (0 => "00111001", 1 => "00111001", 2 => "00111001", 3 => "00111001", 4 => "00000000"),
            58 => (0 => "00111010", 1 => "00111010", 2 => "00111010", 3 => "00111010", 4 => "00000000"),
            59 => (0 => "00111011", 1 => "00111011", 2 => "00111011", 3 => "00111011", 4 => "00000000"),
            60 => (0 => "00111100", 1 => "00111100", 2 => "00111100", 3 => "00111100", 4 => "00000000"),
            61 => (0 => "00111101", 1 => "00111101", 2 => "00111101", 3 => "00111101", 4 => "00000000"),
            62 => (0 => "00111110", 1 => "00111110", 2 => "00111110", 3 => "00111110", 4 => "00000000"),
            63 => (0 => "00111111", 1 => "00111111", 2 => "00111111", 3 => "00111111", 4 => "00000000"),
            64 => (0 => "01000000", 1 => "01000000", 2 => "01000000", 3 => "01000000", 4 => "00000000"),
            65 => (0 => "01000001", 1 => "01000001", 2 => "01000001", 3 => "01000001", 4 => "00000000"),
            66 => (0 => "01000010", 1 => "01000010", 2 => "01000010", 3 => "01000010", 4 => "00000000"),
            67 => (0 => "01000011", 1 => "01000011", 2 => "01000011", 3 => "01000011", 4 => "00000000"),
            68 => (0 => "01000100", 1 => "01000100", 2 => "01000100", 3 => "01000100", 4 => "00000000"),
            69 => (0 => "01000101", 1 => "01000101", 2 => "01000101", 3 => "01000101", 4 => "00000000"),
            70 => (0 => "01000110", 1 => "01000110", 2 => "01000110", 3 => "01000110", 4 => "00000000"),
            71 => (0 => "01000111", 1 => "01000111", 2 => "01000111", 3 => "01000111", 4 => "00000000"),
            72 => (0 => "01001000", 1 => "01001000", 2 => "01001000", 3 => "01001000", 4 => "00000000"),
            73 => (0 => "01001001", 1 => "01001001", 2 => "01001001", 3 => "01001001", 4 => "00000000"),
            74 => (0 => "01001010", 1 => "01001010", 2 => "01001010", 3 => "01001010", 4 => "00000000"),
            75 => (0 => "01001011", 1 => "01001011", 2 => "01001011", 3 => "01001011", 4 => "00000000"),
            76 => (0 => "01001100", 1 => "01001100", 2 => "01001100", 3 => "01001100", 4 => "00000000"),
            77 => (0 => "01001101", 1 => "01001101", 2 => "01001101", 3 => "01001101", 4 => "00000000"),
            78 => (0 => "01001110", 1 => "01001110", 2 => "01001110", 3 => "01001110", 4 => "00000000"),
            79 => (0 => "01001111", 1 => "01001111", 2 => "01001111", 3 => "01001111", 4 => "00000000"),
            80 => (0 => "01010000", 1 => "01010000", 2 => "01010000", 3 => "01010000", 4 => "00000000"),
            81 => (0 => "01010001", 1 => "01010001", 2 => "01010001", 3 => "01010001", 4 => "00000000"),
            82 => (0 => "01010010", 1 => "01010010", 2 => "01010010", 3 => "01010010", 4 => "00000000"),
            83 => (0 => "01010011", 1 => "01010011", 2 => "01010011", 3 => "01010011", 4 => "00000000"),
            84 => (0 => "01010100", 1 => "01010100", 2 => "01010100", 3 => "01010100", 4 => "00000000"),
            85 => (0 => "01010101", 1 => "01010101", 2 => "01010101", 3 => "01010101", 4 => "00000000"),
            86 => (0 => "01010110", 1 => "01010110", 2 => "01010110", 3 => "01010110", 4 => "00000000"),
            87 => (0 => "01010111", 1 => "01010111", 2 => "01010111", 3 => "01010111", 4 => "00000000"),
            88 => (0 => "01011000", 1 => "01011000", 2 => "01011000", 3 => "01011000", 4 => "00000000"),
            89 => (0 => "01011001", 1 => "01011001", 2 => "01011001", 3 => "01011001", 4 => "00000000"),
            90 => (0 => "01011010", 1 => "01011010", 2 => "01011010", 3 => "01011010", 4 => "00000000"),
            91 => (0 => "01011011", 1 => "01011011", 2 => "01011011", 3 => "01011011", 4 => "00000000"),
            92 => (0 => "01011100", 1 => "01011100", 2 => "01011100", 3 => "01011100", 4 => "00000000"),
            93 => (0 => "01011101", 1 => "01011101", 2 => "01011101", 3 => "01011101", 4 => "00000000"),
            94 => (0 => "01011110", 1 => "01011110", 2 => "01011110", 3 => "01011110", 4 => "00000000"),
            95 => (0 => "01011111", 1 => "01011111", 2 => "01011111", 3 => "01011111", 4 => "00000000"),
            96 => (0 => "01100000", 1 => "01100000", 2 => "01100000", 3 => "01100000", 4 => "00000000"),
            97 => (0 => "01100001", 1 => "01100001", 2 => "01100001", 3 => "01100001", 4 => "00000000"),
            98 => (0 => "01100010", 1 => "01100010", 2 => "01100010", 3 => "01100010", 4 => "00000000"),
            99 => (0 => "01100011", 1 => "01100011", 2 => "01100011", 3 => "01100011", 4 => "00000000"),
            100 => (0 => "01100100", 1 => "01100100", 2 => "01100100", 3 => "01100100", 4 => "00000000"),
            101 => (0 => "01100101", 1 => "01100101", 2 => "01100101", 3 => "01100101", 4 => "00000000"),
            102 => (0 => "01100110", 1 => "01100110", 2 => "01100110", 3 => "01100110", 4 => "00000000"),
            103 => (0 => "01100111", 1 => "01100111", 2 => "01100111", 3 => "01100111", 4 => "00000000"),
            104 => (0 => "01101000", 1 => "01101000", 2 => "01101000", 3 => "01101000", 4 => "00000000"),
            105 => (0 => "01101001", 1 => "01101001", 2 => "01101001", 3 => "01101001", 4 => "00000000"),
            106 => (0 => "01101010", 1 => "01101010", 2 => "01101010", 3 => "01101010", 4 => "00000000"),
            107 => (0 => "01101011", 1 => "01101011", 2 => "01101011", 3 => "01101011", 4 => "00000000"),
            108 => (0 => "01101100", 1 => "01101100", 2 => "01101100", 3 => "01101100", 4 => "00000000"),
            109 => (0 => "01101101", 1 => "01101101", 2 => "01101101", 3 => "01101101", 4 => "00000000"),
            110 => (0 => "01101110", 1 => "01101110", 2 => "01101110", 3 => "01101110", 4 => "00000000"),
            111 => (0 => "01101111", 1 => "01101111", 2 => "01101111", 3 => "01101111", 4 => "00000000"),
            112 => (0 => "01110000", 1 => "01110000", 2 => "01110000", 3 => "01110000", 4 => "00000000"),
            113 => (0 => "01110001", 1 => "01110001", 2 => "01110001", 3 => "01110001", 4 => "00000000"),
            114 => (0 => "01110010", 1 => "01110010", 2 => "01110010", 3 => "01110010", 4 => "00000000"),
            115 => (0 => "01110011", 1 => "01110011", 2 => "01110011", 3 => "01110011", 4 => "00000000"),
            116 => (0 => "01110100", 1 => "01110100", 2 => "01110100", 3 => "01110100", 4 => "00000000"),
            117 => (0 => "01110101", 1 => "01110101", 2 => "01110101", 3 => "01110101", 4 => "00000000"),
            118 => (0 => "01110110", 1 => "01110110", 2 => "01110110", 3 => "01110110", 4 => "00000000"),
            119 => (0 => "01110111", 1 => "01110111", 2 => "01110111", 3 => "01110111", 4 => "00000000"),
            120 => (0 => "01111000", 1 => "01111000", 2 => "01111000", 3 => "01111000", 4 => "00000000"),
            121 => (0 => "01111001", 1 => "01111001", 2 => "01111001", 3 => "01111001", 4 => "00000000"),
            122 => (0 => "01111010", 1 => "01111010", 2 => "01111010", 3 => "01111010", 4 => "00000000"),
            123 => (0 => "01111011", 1 => "01111011", 2 => "01111011", 3 => "01111011", 4 => "00000000"),
            124 => (0 => "01111100", 1 => "01111100", 2 => "01111100", 3 => "01111100", 4 => "00000000"),
            125 => (0 => "01111101", 1 => "01111101", 2 => "01111101", 3 => "01111101", 4 => "00000000"),
            126 => (0 => "01111110", 1 => "01111110", 2 => "01111110", 3 => "01111110", 4 => "00000000"),
            127 => (0 => "01111111", 1 => "01111111", 2 => "01111111", 3 => "01111111", 4 => "00000000"),
            128 => (0 => "10000000", 1 => "10000000", 2 => "10000000", 3 => "10000000", 4 => "00000000"),
            129 => (0 => "10000001", 1 => "10000001", 2 => "10000001", 3 => "10000001", 4 => "00000000"),
            130 => (0 => "10000010", 1 => "10000010", 2 => "10000010", 3 => "10000010", 4 => "00000000"),
            131 => (0 => "10000011", 1 => "10000011", 2 => "10000011", 3 => "10000011", 4 => "00000000"),
            132 => (0 => "10000100", 1 => "10000100", 2 => "10000100", 3 => "10000100", 4 => "00000000"),
            133 => (0 => "10000101", 1 => "10000101", 2 => "10000101", 3 => "10000101", 4 => "00000000"),
            134 => (0 => "10000110", 1 => "10000110", 2 => "10000110", 3 => "10000110", 4 => "00000000"),
            135 => (0 => "10000111", 1 => "10000111", 2 => "10000111", 3 => "10000111", 4 => "00000000"),
            136 => (0 => "10001000", 1 => "10001000", 2 => "10001000", 3 => "10001000", 4 => "00000000"),
            137 => (0 => "10001001", 1 => "10001001", 2 => "10001001", 3 => "10001001", 4 => "00000000"),
            138 => (0 => "10001010", 1 => "10001010", 2 => "10001010", 3 => "10001010", 4 => "00000000"),
            139 => (0 => "10001011", 1 => "10001011", 2 => "10001011", 3 => "10001011", 4 => "00000000"),
            140 => (0 => "10001100", 1 => "10001100", 2 => "10001100", 3 => "10001100", 4 => "00000000"),
            141 => (0 => "10001101", 1 => "10001101", 2 => "10001101", 3 => "10001101", 4 => "00000000"),
            142 => (0 => "10001110", 1 => "10001110", 2 => "10001110", 3 => "10001110", 4 => "00000000"),
            143 => (0 => "10001111", 1 => "10001111", 2 => "10001111", 3 => "10001111", 4 => "00000000"),
            144 => (0 => "10010000", 1 => "10010000", 2 => "10010000", 3 => "10010000", 4 => "00000000"),
            145 => (0 => "10010001", 1 => "10010001", 2 => "10010001", 3 => "10010001", 4 => "00000000"),
            146 => (0 => "10010010", 1 => "10010010", 2 => "10010010", 3 => "10010010", 4 => "00000000"),
            147 => (0 => "10010011", 1 => "10010011", 2 => "10010011", 3 => "10010011", 4 => "00000000"),
            148 => (0 => "10010100", 1 => "10010100", 2 => "10010100", 3 => "10010100", 4 => "00000000"),
            149 => (0 => "10010101", 1 => "10010101", 2 => "10010101", 3 => "10010101", 4 => "00000000"),
            150 => (0 => "10010110", 1 => "10010110", 2 => "10010110", 3 => "10010110", 4 => "00000000"),
            151 => (0 => "10010111", 1 => "10010111", 2 => "10010111", 3 => "10010111", 4 => "00000000"),
            152 => (0 => "10011000", 1 => "10011000", 2 => "10011000", 3 => "10011000", 4 => "00000000"),
            153 => (0 => "10011001", 1 => "10011001", 2 => "10011001", 3 => "10011001", 4 => "00000000"),
            154 => (0 => "10011010", 1 => "10011010", 2 => "10011010", 3 => "10011010", 4 => "00000000"),
            155 => (0 => "10011011", 1 => "10011011", 2 => "10011011", 3 => "10011011", 4 => "00000000"),
            156 => (0 => "10011100", 1 => "10011100", 2 => "10011100", 3 => "10011100", 4 => "00000000"),
            157 => (0 => "10011101", 1 => "10011101", 2 => "10011101", 3 => "10011101", 4 => "00000000"),
            158 => (0 => "10011110", 1 => "10011110", 2 => "10011110", 3 => "10011110", 4 => "00000000"),
            159 => (0 => "10011111", 1 => "10011111", 2 => "10011111", 3 => "10011111", 4 => "00000000"),
            160 => (0 => "10100000", 1 => "10100000", 2 => "10100000", 3 => "10100000", 4 => "00000000"),
            161 => (0 => "10100001", 1 => "10100001", 2 => "10100001", 3 => "10100001", 4 => "00000000"),
            162 => (0 => "10100010", 1 => "10100010", 2 => "10100010", 3 => "10100010", 4 => "00000000"),
            163 => (0 => "10100011", 1 => "10100011", 2 => "10100011", 3 => "10100011", 4 => "00000000"),
            164 => (0 => "10100100", 1 => "10100100", 2 => "10100100", 3 => "10100100", 4 => "00000000"),
            165 => (0 => "10100101", 1 => "10100101", 2 => "10100101", 3 => "10100101", 4 => "00000000"),
            166 => (0 => "10100110", 1 => "10100110", 2 => "10100110", 3 => "10100110", 4 => "00000000"),
            167 => (0 => "10100111", 1 => "10100111", 2 => "10100111", 3 => "10100111", 4 => "00000000"),
            168 => (0 => "10101000", 1 => "10101000", 2 => "10101000", 3 => "10101000", 4 => "00000000"),
            169 => (0 => "10101001", 1 => "10101001", 2 => "10101001", 3 => "10101001", 4 => "00000000"),
            170 => (0 => "10101010", 1 => "10101010", 2 => "10101010", 3 => "10101010", 4 => "00000000"),
            171 => (0 => "10101011", 1 => "10101011", 2 => "10101011", 3 => "10101011", 4 => "00000000"),
            172 => (0 => "10101100", 1 => "10101100", 2 => "10101100", 3 => "10101100", 4 => "00000000"),
            173 => (0 => "10101101", 1 => "10101101", 2 => "10101101", 3 => "10101101", 4 => "00000000"),
            174 => (0 => "10101110", 1 => "10101110", 2 => "10101110", 3 => "10101110", 4 => "00000000"),
            175 => (0 => "10101111", 1 => "10101111", 2 => "10101111", 3 => "10101111", 4 => "00000000"),
            176 => (0 => "10110000", 1 => "10110000", 2 => "10110000", 3 => "10110000", 4 => "00000000"),
            177 => (0 => "10110001", 1 => "10110001", 2 => "10110001", 3 => "10110001", 4 => "00000000"),
            178 => (0 => "10110010", 1 => "10110010", 2 => "10110010", 3 => "10110010", 4 => "00000000"),
            179 => (0 => "10110011", 1 => "10110011", 2 => "10110011", 3 => "10110011", 4 => "00000000"),
            180 => (0 => "10110100", 1 => "10110100", 2 => "10110100", 3 => "10110100", 4 => "00000000"),
            181 => (0 => "10110101", 1 => "10110101", 2 => "10110101", 3 => "10110101", 4 => "00000000"),
            182 => (0 => "10110110", 1 => "10110110", 2 => "10110110", 3 => "10110110", 4 => "00000000"),
            183 => (0 => "10110111", 1 => "10110111", 2 => "10110111", 3 => "10110111", 4 => "00000000"),
            184 => (0 => "10111000", 1 => "10111000", 2 => "10111000", 3 => "10111000", 4 => "00000000"),
            185 => (0 => "10111001", 1 => "10111001", 2 => "10111001", 3 => "10111001", 4 => "00000000"),
            186 => (0 => "10111010", 1 => "10111010", 2 => "10111010", 3 => "10111010", 4 => "00000000"),
            187 => (0 => "10111011", 1 => "10111011", 2 => "10111011", 3 => "10111011", 4 => "00000000"),
            188 => (0 => "10111100", 1 => "10111100", 2 => "10111100", 3 => "10111100", 4 => "00000000"),
            189 => (0 => "10111101", 1 => "10111101", 2 => "10111101", 3 => "10111101", 4 => "00000000"),
            190 => (0 => "10111110", 1 => "10111110", 2 => "10111110", 3 => "10111110", 4 => "00000000"),
            191 => (0 => "10111111", 1 => "10111111", 2 => "10111111", 3 => "10111111", 4 => "00000000"),
            192 => (0 => "11000000", 1 => "11000000", 2 => "11000000", 3 => "11000000", 4 => "00000000"),
            193 => (0 => "11000001", 1 => "11000001", 2 => "11000001", 3 => "11000001", 4 => "00000000"),
            194 => (0 => "11000010", 1 => "11000010", 2 => "11000010", 3 => "11000010", 4 => "00000000"),
            195 => (0 => "11000011", 1 => "11000011", 2 => "11000011", 3 => "11000011", 4 => "00000000"),
            196 => (0 => "11000100", 1 => "11000100", 2 => "11000100", 3 => "11000100", 4 => "00000000"),
            197 => (0 => "11000101", 1 => "11000101", 2 => "11000101", 3 => "11000101", 4 => "00000000"),
            198 => (0 => "11000110", 1 => "11000110", 2 => "11000110", 3 => "11000110", 4 => "00000000"),
            199 => (0 => "11000111", 1 => "11000111", 2 => "11000111", 3 => "11000111", 4 => "00000000"),
            200 => (0 => "11001000", 1 => "11001000", 2 => "11001000", 3 => "11001000", 4 => "00000000"),
            201 => (0 => "11001001", 1 => "11001001", 2 => "11001001", 3 => "11001001", 4 => "00000000"),
            202 => (0 => "11001010", 1 => "11001010", 2 => "11001010", 3 => "11001010", 4 => "00000000"),
            203 => (0 => "11001011", 1 => "11001011", 2 => "11001011", 3 => "11001011", 4 => "00000000"),
            204 => (0 => "11001100", 1 => "11001100", 2 => "11001100", 3 => "11001100", 4 => "00000000"),
            205 => (0 => "11001101", 1 => "11001101", 2 => "11001101", 3 => "11001101", 4 => "00000000"),
            206 => (0 => "11001110", 1 => "11001110", 2 => "11001110", 3 => "11001110", 4 => "00000000"),
            207 => (0 => "11001111", 1 => "11001111", 2 => "11001111", 3 => "11001111", 4 => "00000000"),
            208 => (0 => "11010000", 1 => "11010000", 2 => "11010000", 3 => "11010000", 4 => "00000000"),
            209 => (0 => "11010001", 1 => "11010001", 2 => "11010001", 3 => "11010001", 4 => "00000000"),
            210 => (0 => "11010010", 1 => "11010010", 2 => "11010010", 3 => "11010010", 4 => "00000000"),
            211 => (0 => "11010011", 1 => "11010011", 2 => "11010011", 3 => "11010011", 4 => "00000000"),
            212 => (0 => "11010100", 1 => "11010100", 2 => "11010100", 3 => "11010100", 4 => "00000000"),
            213 => (0 => "11010101", 1 => "11010101", 2 => "11010101", 3 => "11010101", 4 => "00000000"),
            214 => (0 => "11010110", 1 => "11010110", 2 => "11010110", 3 => "11010110", 4 => "00000000"),
            215 => (0 => "11010111", 1 => "11010111", 2 => "11010111", 3 => "11010111", 4 => "00000000"),
            216 => (0 => "11011000", 1 => "11011000", 2 => "11011000", 3 => "11011000", 4 => "00000000"),
            217 => (0 => "11011001", 1 => "11011001", 2 => "11011001", 3 => "11011001", 4 => "00000000"),
            218 => (0 => "11011010", 1 => "11011010", 2 => "11011010", 3 => "11011010", 4 => "00000000"),
            219 => (0 => "11011011", 1 => "11011011", 2 => "11011011", 3 => "11011011", 4 => "00000000"),
            220 => (0 => "11011100", 1 => "11011100", 2 => "11011100", 3 => "11011100", 4 => "00000000"),
            221 => (0 => "11011101", 1 => "11011101", 2 => "11011101", 3 => "11011101", 4 => "00000000"),
            222 => (0 => "11011110", 1 => "11011110", 2 => "11011110", 3 => "11011110", 4 => "00000000"),
            223 => (0 => "11011111", 1 => "11011111", 2 => "11011111", 3 => "11011111", 4 => "00000000"),
            224 => (0 => "11100000", 1 => "11100000", 2 => "11100000", 3 => "11100000", 4 => "00000000"),
            225 => (0 => "11100001", 1 => "11100001", 2 => "11100001", 3 => "11100001", 4 => "00000000"),
            226 => (0 => "11100010", 1 => "11100010", 2 => "11100010", 3 => "11100010", 4 => "00000000"),
            227 => (0 => "11100011", 1 => "11100011", 2 => "11100011", 3 => "11100011", 4 => "00000000"),
            228 => (0 => "11100100", 1 => "11100100", 2 => "11100100", 3 => "11100100", 4 => "00000000"),
            229 => (0 => "11100101", 1 => "11100101", 2 => "11100101", 3 => "11100101", 4 => "00000000"),
            230 => (0 => "11100110", 1 => "11100110", 2 => "11100110", 3 => "11100110", 4 => "00000000"),
            231 => (0 => "11100111", 1 => "11100111", 2 => "11100111", 3 => "11100111", 4 => "00000000"),
            232 => (0 => "11101000", 1 => "11101000", 2 => "11101000", 3 => "11101000", 4 => "00000000"),
            233 => (0 => "11101001", 1 => "11101001", 2 => "11101001", 3 => "11101001", 4 => "00000000"),
            234 => (0 => "11101010", 1 => "11101010", 2 => "11101010", 3 => "11101010", 4 => "00000000"),
            235 => (0 => "11101011", 1 => "11101011", 2 => "11101011", 3 => "11101011", 4 => "00000000"),
            236 => (0 => "11101100", 1 => "11101100", 2 => "11101100", 3 => "11101100", 4 => "00000000"),
            237 => (0 => "11101101", 1 => "11101101", 2 => "11101101", 3 => "11101101", 4 => "00000000"),
            238 => (0 => "11101110", 1 => "11101110", 2 => "11101110", 3 => "11101110", 4 => "00000000"),
            239 => (0 => "11101111", 1 => "11101111", 2 => "11101111", 3 => "11101111", 4 => "00000000"),
            240 => (0 => "11110000", 1 => "11110000", 2 => "11110000", 3 => "11110000", 4 => "00000000"),
            241 => (0 => "11110001", 1 => "11110001", 2 => "11110001", 3 => "11110001", 4 => "00000000"),
            242 => (0 => "11110010", 1 => "11110010", 2 => "11110010", 3 => "11110010", 4 => "00000000"),
            243 => (0 => "11110011", 1 => "11110011", 2 => "11110011", 3 => "11110011", 4 => "00000000"),
            244 => (0 => "11110100", 1 => "11110100", 2 => "11110100", 3 => "11110100", 4 => "00000000"),
            245 => (0 => "11110101", 1 => "11110101", 2 => "11110101", 3 => "11110101", 4 => "00000000"),
            246 => (0 => "11110110", 1 => "11110110", 2 => "11110110", 3 => "11110110", 4 => "00000000"),
            247 => (0 => "11110111", 1 => "11110111", 2 => "11110111", 3 => "11110111", 4 => "00000000"),
            248 => (0 => "11111000", 1 => "11111000", 2 => "11111000", 3 => "11111000", 4 => "00000000"),
            249 => (0 => "11111001", 1 => "11111001", 2 => "11111001", 3 => "11111001", 4 => "00000000"),
            250 => (0 => "11111010", 1 => "11111010", 2 => "11111010", 3 => "11111010", 4 => "00000000"),
            251 => (0 => "11111011", 1 => "11111011", 2 => "11111011", 3 => "11111011", 4 => "00000000"),
            252 => (0 => "11111100", 1 => "11111100", 2 => "11111100", 3 => "11111100", 4 => "00000000"),
            253 => (0 => "11111101", 1 => "11111101", 2 => "11111101", 3 => "11111101", 4 => "00000000"),
            254 => (0 => "11111110", 1 => "11111110", 2 => "11111110", 3 => "11111110", 4 => "00000000"),
            255 => (0 => "11111111", 1 => "11111111", 2 => "11111111", 3 => "11111111", 4 => "00000000")
    );
	
	-- 0 => "00000000" & "000"  & "0000",
	constant output : outputvect_t := (
	                0 => "000000000000000",
            1 => "000000010000111",
            2 => "000000100001001",
            3 => "000000110001110",
            4 => "000001000001010",
            5 => "000001010001101",
            6 => "000001100000011",
            7 => "000001110000100",
            8 => "000010000001011",
            9 => "000010010001100",
            10 => "000010100000010",
            11 => "000010110000101",
            12 => "000011000000001",
            13 => "000011010000110",
            14 => "000011100001000",
            15 => "000011110001111",
            16 => "000100000001100",
            17 => "000100010001011",
            18 => "000100100000101",
            19 => "000100110000010",
            20 => "000101000000110",
            21 => "000101010000001",
            22 => "000101100001111",
            23 => "000101110001000",
            24 => "000110000000111",
            25 => "000110010000000",
            26 => "000110100001110",
            27 => "000110110001001",
            28 => "000111000001101",
            29 => "000111010001010",
            30 => "000111100000100",
            31 => "000111110000011",
            32 => "001000000001101",
            33 => "001000010001010",
            34 => "001000100000100",
            35 => "001000110000011",
            36 => "001001000000111",
            37 => "001001010000000",
            38 => "001001100001110",
            39 => "001001110001001",
            40 => "001010000000110",
            41 => "001010010000001",
            42 => "001010100001111",
            43 => "001010110001000",
            44 => "001011000001100",
            45 => "001011010001011",
            46 => "001011100000101",
            47 => "001011110000010",
            48 => "001100000000001",
            49 => "001100010000110",
            50 => "001100100001000",
            51 => "001100110001111",
            52 => "001101000001011",
            53 => "001101010001100",
            54 => "001101100000010",
            55 => "001101110000101",
            56 => "001110000001010",
            57 => "001110010001101",
            58 => "001110100000011",
            59 => "001110110000100",
            60 => "001111000000000",
            61 => "001111010000111",
            62 => "001111100001001",
            63 => "001111110001110",
            64 => "010000000001110",
            65 => "010000010001001",
            66 => "010000100000111",
            67 => "010000110000000",
            68 => "010001000000100",
            69 => "010001010000011",
            70 => "010001100001101",
            71 => "010001110001010",
            72 => "010010000000101",
            73 => "010010010000010",
            74 => "010010100001100",
            75 => "010010110001011",
            76 => "010011000001111",
            77 => "010011010001000",
            78 => "010011100000110",
            79 => "010011110000001",
            80 => "010100000000010",
            81 => "010100010000101",
            82 => "010100100001011",
            83 => "010100110001100",
            84 => "010101000001000",
            85 => "010101010001111",
            86 => "010101100000001",
            87 => "010101110000110",
            88 => "010110000001001",
            89 => "010110010001110",
            90 => "010110100000000",
            91 => "010110110000111",
            92 => "010111000000011",
            93 => "010111010000100",
            94 => "010111100001010",
            95 => "010111110001101",
            96 => "011000000000011",
            97 => "011000010000100",
            98 => "011000100001010",
            99 => "011000110001101",
            100 => "011001000001001",
            101 => "011001010001110",
            102 => "011001100000000",
            103 => "011001110000111",
            104 => "011010000001000",
            105 => "011010010001111",
            106 => "011010100000001",
            107 => "011010110000110",
            108 => "011011000000010",
            109 => "011011010000101",
            110 => "011011100001011",
            111 => "011011110001100",
            112 => "011100000001111",
            113 => "011100010001000",
            114 => "011100100000110",
            115 => "011100110000001",
            116 => "011101000000101",
            117 => "011101010000010",
            118 => "011101100001100",
            119 => "011101110001011",
            120 => "011110000000100",
            121 => "011110010000011",
            122 => "011110100001101",
            123 => "011110110001010",
            124 => "011111000001110",
            125 => "011111010001001",
            126 => "011111100000111",
            127 => "011111110000000",
            128 => "100000000001111",
            129 => "100000010001000",
            130 => "100000100000110",
            131 => "100000110000001",
            132 => "100001000000101",
            133 => "100001010000010",
            134 => "100001100001100",
            135 => "100001110001011",
            136 => "100010000000100",
            137 => "100010010000011",
            138 => "100010100001101",
            139 => "100010110001010",
            140 => "100011000001110",
            141 => "100011010001001",
            142 => "100011100000111",
            143 => "100011110000000",
            144 => "100100000000011",
            145 => "100100010000100",
            146 => "100100100001010",
            147 => "100100110001101",
            148 => "100101000001001",
            149 => "100101010001110",
            150 => "100101100000000",
            151 => "100101110000111",
            152 => "100110000001000",
            153 => "100110010001111",
            154 => "100110100000001",
            155 => "100110110000110",
            156 => "100111000000010",
            157 => "100111010000101",
            158 => "100111100001011",
            159 => "100111110001100",
            160 => "101000000000010",
            161 => "101000010000101",
            162 => "101000100001011",
            163 => "101000110001100",
            164 => "101001000001000",
            165 => "101001010001111",
            166 => "101001100000001",
            167 => "101001110000110",
            168 => "101010000001001",
            169 => "101010010001110",
            170 => "101010100000000",
            171 => "101010110000111",
            172 => "101011000000011",
            173 => "101011010000100",
            174 => "101011100001010",
            175 => "101011110001101",
            176 => "101100000001110",
            177 => "101100010001001",
            178 => "101100100000111",
            179 => "101100110000000",
            180 => "101101000000100",
            181 => "101101010000011",
            182 => "101101100001101",
            183 => "101101110001010",
            184 => "101110000000101",
            185 => "101110010000010",
            186 => "101110100001100",
            187 => "101110110001011",
            188 => "101111000001111",
            189 => "101111010001000",
            190 => "101111100000110",
            191 => "101111110000001",
            192 => "110000000000001",
            193 => "110000010000110",
            194 => "110000100001000",
            195 => "110000110001111",
            196 => "110001000001011",
            197 => "110001010001100",
            198 => "110001100000010",
            199 => "110001110000101",
            200 => "110010000001010",
            201 => "110010010001101",
            202 => "110010100000011",
            203 => "110010110000100",
            204 => "110011000000000",
            205 => "110011010000111",
            206 => "110011100001001",
            207 => "110011110001110",
            208 => "110100000001101",
            209 => "110100010001010",
            210 => "110100100000100",
            211 => "110100110000011",
            212 => "110101000000111",
            213 => "110101010000000",
            214 => "110101100001110",
            215 => "110101110001001",
            216 => "110110000000110",
            217 => "110110010000001",
            218 => "110110100001111",
            219 => "110110110001000",
            220 => "110111000001100",
            221 => "110111010001011",
            222 => "110111100000101",
            223 => "110111110000010",
            224 => "111000000001100",
            225 => "111000010001011",
            226 => "111000100000101",
            227 => "111000110000010",
            228 => "111001000000110",
            229 => "111001010000001",
            230 => "111001100001111",
            231 => "111001110001000",
            232 => "111010000000111",
            233 => "111010010000000",
            234 => "111010100001110",
            235 => "111010110001001",
            236 => "111011000001101",
            237 => "111011010001010",
            238 => "111011100000100",
            239 => "111011110000011",
            240 => "111100000000000",
            241 => "111100010000111",
            242 => "111100100001001",
            243 => "111100110001110",
            244 => "111101000001010",
            245 => "111101010001101",
            246 => "111101100000011",
            247 => "111101110000100",
            248 => "111110000001011",
            249 => "111110010001100",
            250 => "111110100000010",
            251 => "111110110000101",
            252 => "111111000000001",
            253 => "111111010000110",
            254 => "111111100001000",
            255 => "111111110001111"
	);
end package;
