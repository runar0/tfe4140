library ieee;
use ieee.std_logic_1164.all;

package liaison_tb_data is

    constant count : integer := 4096;

    type inputvect_t is array(0 to count-1, 0 to 4) of std_logic_vector(7 downto 0);
    type outputvect_t is array(0 to count-1) of std_logic_vector(14 downto 0);

    -- 0 => (0 => "00000000", 1 => "00000000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
    constant input : inputvect_t := (
                    0 => (0 => "00000000", 1 => "00000000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            1 => (0 => "00000001", 1 => "00000001", 2 => "00000001", 3 => "00000001", 4 => "00000000"),
            2 => (0 => "00000010", 1 => "00000010", 2 => "00000010", 3 => "00000010", 4 => "00000000"),
            3 => (0 => "00000011", 1 => "00000011", 2 => "00000011", 3 => "00000011", 4 => "00000000"),
            4 => (0 => "00000100", 1 => "00000100", 2 => "00000100", 3 => "00000100", 4 => "00000000"),
            5 => (0 => "00000101", 1 => "00000101", 2 => "00000101", 3 => "00000101", 4 => "00000000"),
            6 => (0 => "00000110", 1 => "00000110", 2 => "00000110", 3 => "00000110", 4 => "00000000"),
            7 => (0 => "00000111", 1 => "00000111", 2 => "00000111", 3 => "00000111", 4 => "00000000"),
            8 => (0 => "00001000", 1 => "00001000", 2 => "00001000", 3 => "00001000", 4 => "00000000"),
            9 => (0 => "00001001", 1 => "00001001", 2 => "00001001", 3 => "00001001", 4 => "00000000"),
            10 => (0 => "00001010", 1 => "00001010", 2 => "00001010", 3 => "00001010", 4 => "00000000"),
            11 => (0 => "00001011", 1 => "00001011", 2 => "00001011", 3 => "00001011", 4 => "00000000"),
            12 => (0 => "00001100", 1 => "00001100", 2 => "00001100", 3 => "00001100", 4 => "00000000"),
            13 => (0 => "00001101", 1 => "00001101", 2 => "00001101", 3 => "00001101", 4 => "00000000"),
            14 => (0 => "00001110", 1 => "00001110", 2 => "00001110", 3 => "00001110", 4 => "00000000"),
            15 => (0 => "00001111", 1 => "00001111", 2 => "00001111", 3 => "00001111", 4 => "00000000"),
            16 => (0 => "00010000", 1 => "00010000", 2 => "00010000", 3 => "00010000", 4 => "00000000"),
            17 => (0 => "00010001", 1 => "00010001", 2 => "00010001", 3 => "00010001", 4 => "00000000"),
            18 => (0 => "00010010", 1 => "00010010", 2 => "00010010", 3 => "00010010", 4 => "00000000"),
            19 => (0 => "00010011", 1 => "00010011", 2 => "00010011", 3 => "00010011", 4 => "00000000"),
            20 => (0 => "00010100", 1 => "00010100", 2 => "00010100", 3 => "00010100", 4 => "00000000"),
            21 => (0 => "00010101", 1 => "00010101", 2 => "00010101", 3 => "00010101", 4 => "00000000"),
            22 => (0 => "00010110", 1 => "00010110", 2 => "00010110", 3 => "00010110", 4 => "00000000"),
            23 => (0 => "00010111", 1 => "00010111", 2 => "00010111", 3 => "00010111", 4 => "00000000"),
            24 => (0 => "00011000", 1 => "00011000", 2 => "00011000", 3 => "00011000", 4 => "00000000"),
            25 => (0 => "00011001", 1 => "00011001", 2 => "00011001", 3 => "00011001", 4 => "00000000"),
            26 => (0 => "00011010", 1 => "00011010", 2 => "00011010", 3 => "00011010", 4 => "00000000"),
            27 => (0 => "00011011", 1 => "00011011", 2 => "00011011", 3 => "00011011", 4 => "00000000"),
            28 => (0 => "00011100", 1 => "00011100", 2 => "00011100", 3 => "00011100", 4 => "00000000"),
            29 => (0 => "00011101", 1 => "00011101", 2 => "00011101", 3 => "00011101", 4 => "00000000"),
            30 => (0 => "00011110", 1 => "00011110", 2 => "00011110", 3 => "00011110", 4 => "00000000"),
            31 => (0 => "00011111", 1 => "00011111", 2 => "00011111", 3 => "00011111", 4 => "00000000"),
            32 => (0 => "00100000", 1 => "00100000", 2 => "00100000", 3 => "00100000", 4 => "00000000"),
            33 => (0 => "00100001", 1 => "00100001", 2 => "00100001", 3 => "00100001", 4 => "00000000"),
            34 => (0 => "00100010", 1 => "00100010", 2 => "00100010", 3 => "00100010", 4 => "00000000"),
            35 => (0 => "00100011", 1 => "00100011", 2 => "00100011", 3 => "00100011", 4 => "00000000"),
            36 => (0 => "00100100", 1 => "00100100", 2 => "00100100", 3 => "00100100", 4 => "00000000"),
            37 => (0 => "00100101", 1 => "00100101", 2 => "00100101", 3 => "00100101", 4 => "00000000"),
            38 => (0 => "00100110", 1 => "00100110", 2 => "00100110", 3 => "00100110", 4 => "00000000"),
            39 => (0 => "00100111", 1 => "00100111", 2 => "00100111", 3 => "00100111", 4 => "00000000"),
            40 => (0 => "00101000", 1 => "00101000", 2 => "00101000", 3 => "00101000", 4 => "00000000"),
            41 => (0 => "00101001", 1 => "00101001", 2 => "00101001", 3 => "00101001", 4 => "00000000"),
            42 => (0 => "00101010", 1 => "00101010", 2 => "00101010", 3 => "00101010", 4 => "00000000"),
            43 => (0 => "00101011", 1 => "00101011", 2 => "00101011", 3 => "00101011", 4 => "00000000"),
            44 => (0 => "00101100", 1 => "00101100", 2 => "00101100", 3 => "00101100", 4 => "00000000"),
            45 => (0 => "00101101", 1 => "00101101", 2 => "00101101", 3 => "00101101", 4 => "00000000"),
            46 => (0 => "00101110", 1 => "00101110", 2 => "00101110", 3 => "00101110", 4 => "00000000"),
            47 => (0 => "00101111", 1 => "00101111", 2 => "00101111", 3 => "00101111", 4 => "00000000"),
            48 => (0 => "00110000", 1 => "00110000", 2 => "00110000", 3 => "00110000", 4 => "00000000"),
            49 => (0 => "00110001", 1 => "00110001", 2 => "00110001", 3 => "00110001", 4 => "00000000"),
            50 => (0 => "00110010", 1 => "00110010", 2 => "00110010", 3 => "00110010", 4 => "00000000"),
            51 => (0 => "00110011", 1 => "00110011", 2 => "00110011", 3 => "00110011", 4 => "00000000"),
            52 => (0 => "00110100", 1 => "00110100", 2 => "00110100", 3 => "00110100", 4 => "00000000"),
            53 => (0 => "00110101", 1 => "00110101", 2 => "00110101", 3 => "00110101", 4 => "00000000"),
            54 => (0 => "00110110", 1 => "00110110", 2 => "00110110", 3 => "00110110", 4 => "00000000"),
            55 => (0 => "00110111", 1 => "00110111", 2 => "00110111", 3 => "00110111", 4 => "00000000"),
            56 => (0 => "00111000", 1 => "00111000", 2 => "00111000", 3 => "00111000", 4 => "00000000"),
            57 => (0 => "00111001", 1 => "00111001", 2 => "00111001", 3 => "00111001", 4 => "00000000"),
            58 => (0 => "00111010", 1 => "00111010", 2 => "00111010", 3 => "00111010", 4 => "00000000"),
            59 => (0 => "00111011", 1 => "00111011", 2 => "00111011", 3 => "00111011", 4 => "00000000"),
            60 => (0 => "00111100", 1 => "00111100", 2 => "00111100", 3 => "00111100", 4 => "00000000"),
            61 => (0 => "00111101", 1 => "00111101", 2 => "00111101", 3 => "00111101", 4 => "00000000"),
            62 => (0 => "00111110", 1 => "00111110", 2 => "00111110", 3 => "00111110", 4 => "00000000"),
            63 => (0 => "00111111", 1 => "00111111", 2 => "00111111", 3 => "00111111", 4 => "00000000"),
            64 => (0 => "01000000", 1 => "01000000", 2 => "01000000", 3 => "01000000", 4 => "00000000"),
            65 => (0 => "01000001", 1 => "01000001", 2 => "01000001", 3 => "01000001", 4 => "00000000"),
            66 => (0 => "01000010", 1 => "01000010", 2 => "01000010", 3 => "01000010", 4 => "00000000"),
            67 => (0 => "01000011", 1 => "01000011", 2 => "01000011", 3 => "01000011", 4 => "00000000"),
            68 => (0 => "01000100", 1 => "01000100", 2 => "01000100", 3 => "01000100", 4 => "00000000"),
            69 => (0 => "01000101", 1 => "01000101", 2 => "01000101", 3 => "01000101", 4 => "00000000"),
            70 => (0 => "01000110", 1 => "01000110", 2 => "01000110", 3 => "01000110", 4 => "00000000"),
            71 => (0 => "01000111", 1 => "01000111", 2 => "01000111", 3 => "01000111", 4 => "00000000"),
            72 => (0 => "01001000", 1 => "01001000", 2 => "01001000", 3 => "01001000", 4 => "00000000"),
            73 => (0 => "01001001", 1 => "01001001", 2 => "01001001", 3 => "01001001", 4 => "00000000"),
            74 => (0 => "01001010", 1 => "01001010", 2 => "01001010", 3 => "01001010", 4 => "00000000"),
            75 => (0 => "01001011", 1 => "01001011", 2 => "01001011", 3 => "01001011", 4 => "00000000"),
            76 => (0 => "01001100", 1 => "01001100", 2 => "01001100", 3 => "01001100", 4 => "00000000"),
            77 => (0 => "01001101", 1 => "01001101", 2 => "01001101", 3 => "01001101", 4 => "00000000"),
            78 => (0 => "01001110", 1 => "01001110", 2 => "01001110", 3 => "01001110", 4 => "00000000"),
            79 => (0 => "01001111", 1 => "01001111", 2 => "01001111", 3 => "01001111", 4 => "00000000"),
            80 => (0 => "01010000", 1 => "01010000", 2 => "01010000", 3 => "01010000", 4 => "00000000"),
            81 => (0 => "01010001", 1 => "01010001", 2 => "01010001", 3 => "01010001", 4 => "00000000"),
            82 => (0 => "01010010", 1 => "01010010", 2 => "01010010", 3 => "01010010", 4 => "00000000"),
            83 => (0 => "01010011", 1 => "01010011", 2 => "01010011", 3 => "01010011", 4 => "00000000"),
            84 => (0 => "01010100", 1 => "01010100", 2 => "01010100", 3 => "01010100", 4 => "00000000"),
            85 => (0 => "01010101", 1 => "01010101", 2 => "01010101", 3 => "01010101", 4 => "00000000"),
            86 => (0 => "01010110", 1 => "01010110", 2 => "01010110", 3 => "01010110", 4 => "00000000"),
            87 => (0 => "01010111", 1 => "01010111", 2 => "01010111", 3 => "01010111", 4 => "00000000"),
            88 => (0 => "01011000", 1 => "01011000", 2 => "01011000", 3 => "01011000", 4 => "00000000"),
            89 => (0 => "01011001", 1 => "01011001", 2 => "01011001", 3 => "01011001", 4 => "00000000"),
            90 => (0 => "01011010", 1 => "01011010", 2 => "01011010", 3 => "01011010", 4 => "00000000"),
            91 => (0 => "01011011", 1 => "01011011", 2 => "01011011", 3 => "01011011", 4 => "00000000"),
            92 => (0 => "01011100", 1 => "01011100", 2 => "01011100", 3 => "01011100", 4 => "00000000"),
            93 => (0 => "01011101", 1 => "01011101", 2 => "01011101", 3 => "01011101", 4 => "00000000"),
            94 => (0 => "01011110", 1 => "01011110", 2 => "01011110", 3 => "01011110", 4 => "00000000"),
            95 => (0 => "01011111", 1 => "01011111", 2 => "01011111", 3 => "01011111", 4 => "00000000"),
            96 => (0 => "01100000", 1 => "01100000", 2 => "01100000", 3 => "01100000", 4 => "00000000"),
            97 => (0 => "01100001", 1 => "01100001", 2 => "01100001", 3 => "01100001", 4 => "00000000"),
            98 => (0 => "01100010", 1 => "01100010", 2 => "01100010", 3 => "01100010", 4 => "00000000"),
            99 => (0 => "01100011", 1 => "01100011", 2 => "01100011", 3 => "01100011", 4 => "00000000"),
            100 => (0 => "01100100", 1 => "01100100", 2 => "01100100", 3 => "01100100", 4 => "00000000"),
            101 => (0 => "01100101", 1 => "01100101", 2 => "01100101", 3 => "01100101", 4 => "00000000"),
            102 => (0 => "01100110", 1 => "01100110", 2 => "01100110", 3 => "01100110", 4 => "00000000"),
            103 => (0 => "01100111", 1 => "01100111", 2 => "01100111", 3 => "01100111", 4 => "00000000"),
            104 => (0 => "01101000", 1 => "01101000", 2 => "01101000", 3 => "01101000", 4 => "00000000"),
            105 => (0 => "01101001", 1 => "01101001", 2 => "01101001", 3 => "01101001", 4 => "00000000"),
            106 => (0 => "01101010", 1 => "01101010", 2 => "01101010", 3 => "01101010", 4 => "00000000"),
            107 => (0 => "01101011", 1 => "01101011", 2 => "01101011", 3 => "01101011", 4 => "00000000"),
            108 => (0 => "01101100", 1 => "01101100", 2 => "01101100", 3 => "01101100", 4 => "00000000"),
            109 => (0 => "01101101", 1 => "01101101", 2 => "01101101", 3 => "01101101", 4 => "00000000"),
            110 => (0 => "01101110", 1 => "01101110", 2 => "01101110", 3 => "01101110", 4 => "00000000"),
            111 => (0 => "01101111", 1 => "01101111", 2 => "01101111", 3 => "01101111", 4 => "00000000"),
            112 => (0 => "01110000", 1 => "01110000", 2 => "01110000", 3 => "01110000", 4 => "00000000"),
            113 => (0 => "01110001", 1 => "01110001", 2 => "01110001", 3 => "01110001", 4 => "00000000"),
            114 => (0 => "01110010", 1 => "01110010", 2 => "01110010", 3 => "01110010", 4 => "00000000"),
            115 => (0 => "01110011", 1 => "01110011", 2 => "01110011", 3 => "01110011", 4 => "00000000"),
            116 => (0 => "01110100", 1 => "01110100", 2 => "01110100", 3 => "01110100", 4 => "00000000"),
            117 => (0 => "01110101", 1 => "01110101", 2 => "01110101", 3 => "01110101", 4 => "00000000"),
            118 => (0 => "01110110", 1 => "01110110", 2 => "01110110", 3 => "01110110", 4 => "00000000"),
            119 => (0 => "01110111", 1 => "01110111", 2 => "01110111", 3 => "01110111", 4 => "00000000"),
            120 => (0 => "01111000", 1 => "01111000", 2 => "01111000", 3 => "01111000", 4 => "00000000"),
            121 => (0 => "01111001", 1 => "01111001", 2 => "01111001", 3 => "01111001", 4 => "00000000"),
            122 => (0 => "01111010", 1 => "01111010", 2 => "01111010", 3 => "01111010", 4 => "00000000"),
            123 => (0 => "01111011", 1 => "01111011", 2 => "01111011", 3 => "01111011", 4 => "00000000"),
            124 => (0 => "01111100", 1 => "01111100", 2 => "01111100", 3 => "01111100", 4 => "00000000"),
            125 => (0 => "01111101", 1 => "01111101", 2 => "01111101", 3 => "01111101", 4 => "00000000"),
            126 => (0 => "01111110", 1 => "01111110", 2 => "01111110", 3 => "01111110", 4 => "00000000"),
            127 => (0 => "01111111", 1 => "01111111", 2 => "01111111", 3 => "01111111", 4 => "00000000"),
            128 => (0 => "10000000", 1 => "10000000", 2 => "10000000", 3 => "10000000", 4 => "00000000"),
            129 => (0 => "10000001", 1 => "10000001", 2 => "10000001", 3 => "10000001", 4 => "00000000"),
            130 => (0 => "10000010", 1 => "10000010", 2 => "10000010", 3 => "10000010", 4 => "00000000"),
            131 => (0 => "10000011", 1 => "10000011", 2 => "10000011", 3 => "10000011", 4 => "00000000"),
            132 => (0 => "10000100", 1 => "10000100", 2 => "10000100", 3 => "10000100", 4 => "00000000"),
            133 => (0 => "10000101", 1 => "10000101", 2 => "10000101", 3 => "10000101", 4 => "00000000"),
            134 => (0 => "10000110", 1 => "10000110", 2 => "10000110", 3 => "10000110", 4 => "00000000"),
            135 => (0 => "10000111", 1 => "10000111", 2 => "10000111", 3 => "10000111", 4 => "00000000"),
            136 => (0 => "10001000", 1 => "10001000", 2 => "10001000", 3 => "10001000", 4 => "00000000"),
            137 => (0 => "10001001", 1 => "10001001", 2 => "10001001", 3 => "10001001", 4 => "00000000"),
            138 => (0 => "10001010", 1 => "10001010", 2 => "10001010", 3 => "10001010", 4 => "00000000"),
            139 => (0 => "10001011", 1 => "10001011", 2 => "10001011", 3 => "10001011", 4 => "00000000"),
            140 => (0 => "10001100", 1 => "10001100", 2 => "10001100", 3 => "10001100", 4 => "00000000"),
            141 => (0 => "10001101", 1 => "10001101", 2 => "10001101", 3 => "10001101", 4 => "00000000"),
            142 => (0 => "10001110", 1 => "10001110", 2 => "10001110", 3 => "10001110", 4 => "00000000"),
            143 => (0 => "10001111", 1 => "10001111", 2 => "10001111", 3 => "10001111", 4 => "00000000"),
            144 => (0 => "10010000", 1 => "10010000", 2 => "10010000", 3 => "10010000", 4 => "00000000"),
            145 => (0 => "10010001", 1 => "10010001", 2 => "10010001", 3 => "10010001", 4 => "00000000"),
            146 => (0 => "10010010", 1 => "10010010", 2 => "10010010", 3 => "10010010", 4 => "00000000"),
            147 => (0 => "10010011", 1 => "10010011", 2 => "10010011", 3 => "10010011", 4 => "00000000"),
            148 => (0 => "10010100", 1 => "10010100", 2 => "10010100", 3 => "10010100", 4 => "00000000"),
            149 => (0 => "10010101", 1 => "10010101", 2 => "10010101", 3 => "10010101", 4 => "00000000"),
            150 => (0 => "10010110", 1 => "10010110", 2 => "10010110", 3 => "10010110", 4 => "00000000"),
            151 => (0 => "10010111", 1 => "10010111", 2 => "10010111", 3 => "10010111", 4 => "00000000"),
            152 => (0 => "10011000", 1 => "10011000", 2 => "10011000", 3 => "10011000", 4 => "00000000"),
            153 => (0 => "10011001", 1 => "10011001", 2 => "10011001", 3 => "10011001", 4 => "00000000"),
            154 => (0 => "10011010", 1 => "10011010", 2 => "10011010", 3 => "10011010", 4 => "00000000"),
            155 => (0 => "10011011", 1 => "10011011", 2 => "10011011", 3 => "10011011", 4 => "00000000"),
            156 => (0 => "10011100", 1 => "10011100", 2 => "10011100", 3 => "10011100", 4 => "00000000"),
            157 => (0 => "10011101", 1 => "10011101", 2 => "10011101", 3 => "10011101", 4 => "00000000"),
            158 => (0 => "10011110", 1 => "10011110", 2 => "10011110", 3 => "10011110", 4 => "00000000"),
            159 => (0 => "10011111", 1 => "10011111", 2 => "10011111", 3 => "10011111", 4 => "00000000"),
            160 => (0 => "10100000", 1 => "10100000", 2 => "10100000", 3 => "10100000", 4 => "00000000"),
            161 => (0 => "10100001", 1 => "10100001", 2 => "10100001", 3 => "10100001", 4 => "00000000"),
            162 => (0 => "10100010", 1 => "10100010", 2 => "10100010", 3 => "10100010", 4 => "00000000"),
            163 => (0 => "10100011", 1 => "10100011", 2 => "10100011", 3 => "10100011", 4 => "00000000"),
            164 => (0 => "10100100", 1 => "10100100", 2 => "10100100", 3 => "10100100", 4 => "00000000"),
            165 => (0 => "10100101", 1 => "10100101", 2 => "10100101", 3 => "10100101", 4 => "00000000"),
            166 => (0 => "10100110", 1 => "10100110", 2 => "10100110", 3 => "10100110", 4 => "00000000"),
            167 => (0 => "10100111", 1 => "10100111", 2 => "10100111", 3 => "10100111", 4 => "00000000"),
            168 => (0 => "10101000", 1 => "10101000", 2 => "10101000", 3 => "10101000", 4 => "00000000"),
            169 => (0 => "10101001", 1 => "10101001", 2 => "10101001", 3 => "10101001", 4 => "00000000"),
            170 => (0 => "10101010", 1 => "10101010", 2 => "10101010", 3 => "10101010", 4 => "00000000"),
            171 => (0 => "10101011", 1 => "10101011", 2 => "10101011", 3 => "10101011", 4 => "00000000"),
            172 => (0 => "10101100", 1 => "10101100", 2 => "10101100", 3 => "10101100", 4 => "00000000"),
            173 => (0 => "10101101", 1 => "10101101", 2 => "10101101", 3 => "10101101", 4 => "00000000"),
            174 => (0 => "10101110", 1 => "10101110", 2 => "10101110", 3 => "10101110", 4 => "00000000"),
            175 => (0 => "10101111", 1 => "10101111", 2 => "10101111", 3 => "10101111", 4 => "00000000"),
            176 => (0 => "10110000", 1 => "10110000", 2 => "10110000", 3 => "10110000", 4 => "00000000"),
            177 => (0 => "10110001", 1 => "10110001", 2 => "10110001", 3 => "10110001", 4 => "00000000"),
            178 => (0 => "10110010", 1 => "10110010", 2 => "10110010", 3 => "10110010", 4 => "00000000"),
            179 => (0 => "10110011", 1 => "10110011", 2 => "10110011", 3 => "10110011", 4 => "00000000"),
            180 => (0 => "10110100", 1 => "10110100", 2 => "10110100", 3 => "10110100", 4 => "00000000"),
            181 => (0 => "10110101", 1 => "10110101", 2 => "10110101", 3 => "10110101", 4 => "00000000"),
            182 => (0 => "10110110", 1 => "10110110", 2 => "10110110", 3 => "10110110", 4 => "00000000"),
            183 => (0 => "10110111", 1 => "10110111", 2 => "10110111", 3 => "10110111", 4 => "00000000"),
            184 => (0 => "10111000", 1 => "10111000", 2 => "10111000", 3 => "10111000", 4 => "00000000"),
            185 => (0 => "10111001", 1 => "10111001", 2 => "10111001", 3 => "10111001", 4 => "00000000"),
            186 => (0 => "10111010", 1 => "10111010", 2 => "10111010", 3 => "10111010", 4 => "00000000"),
            187 => (0 => "10111011", 1 => "10111011", 2 => "10111011", 3 => "10111011", 4 => "00000000"),
            188 => (0 => "10111100", 1 => "10111100", 2 => "10111100", 3 => "10111100", 4 => "00000000"),
            189 => (0 => "10111101", 1 => "10111101", 2 => "10111101", 3 => "10111101", 4 => "00000000"),
            190 => (0 => "10111110", 1 => "10111110", 2 => "10111110", 3 => "10111110", 4 => "00000000"),
            191 => (0 => "10111111", 1 => "10111111", 2 => "10111111", 3 => "10111111", 4 => "00000000"),
            192 => (0 => "11000000", 1 => "11000000", 2 => "11000000", 3 => "11000000", 4 => "00000000"),
            193 => (0 => "11000001", 1 => "11000001", 2 => "11000001", 3 => "11000001", 4 => "00000000"),
            194 => (0 => "11000010", 1 => "11000010", 2 => "11000010", 3 => "11000010", 4 => "00000000"),
            195 => (0 => "11000011", 1 => "11000011", 2 => "11000011", 3 => "11000011", 4 => "00000000"),
            196 => (0 => "11000100", 1 => "11000100", 2 => "11000100", 3 => "11000100", 4 => "00000000"),
            197 => (0 => "11000101", 1 => "11000101", 2 => "11000101", 3 => "11000101", 4 => "00000000"),
            198 => (0 => "11000110", 1 => "11000110", 2 => "11000110", 3 => "11000110", 4 => "00000000"),
            199 => (0 => "11000111", 1 => "11000111", 2 => "11000111", 3 => "11000111", 4 => "00000000"),
            200 => (0 => "11001000", 1 => "11001000", 2 => "11001000", 3 => "11001000", 4 => "00000000"),
            201 => (0 => "11001001", 1 => "11001001", 2 => "11001001", 3 => "11001001", 4 => "00000000"),
            202 => (0 => "11001010", 1 => "11001010", 2 => "11001010", 3 => "11001010", 4 => "00000000"),
            203 => (0 => "11001011", 1 => "11001011", 2 => "11001011", 3 => "11001011", 4 => "00000000"),
            204 => (0 => "11001100", 1 => "11001100", 2 => "11001100", 3 => "11001100", 4 => "00000000"),
            205 => (0 => "11001101", 1 => "11001101", 2 => "11001101", 3 => "11001101", 4 => "00000000"),
            206 => (0 => "11001110", 1 => "11001110", 2 => "11001110", 3 => "11001110", 4 => "00000000"),
            207 => (0 => "11001111", 1 => "11001111", 2 => "11001111", 3 => "11001111", 4 => "00000000"),
            208 => (0 => "11010000", 1 => "11010000", 2 => "11010000", 3 => "11010000", 4 => "00000000"),
            209 => (0 => "11010001", 1 => "11010001", 2 => "11010001", 3 => "11010001", 4 => "00000000"),
            210 => (0 => "11010010", 1 => "11010010", 2 => "11010010", 3 => "11010010", 4 => "00000000"),
            211 => (0 => "11010011", 1 => "11010011", 2 => "11010011", 3 => "11010011", 4 => "00000000"),
            212 => (0 => "11010100", 1 => "11010100", 2 => "11010100", 3 => "11010100", 4 => "00000000"),
            213 => (0 => "11010101", 1 => "11010101", 2 => "11010101", 3 => "11010101", 4 => "00000000"),
            214 => (0 => "11010110", 1 => "11010110", 2 => "11010110", 3 => "11010110", 4 => "00000000"),
            215 => (0 => "11010111", 1 => "11010111", 2 => "11010111", 3 => "11010111", 4 => "00000000"),
            216 => (0 => "11011000", 1 => "11011000", 2 => "11011000", 3 => "11011000", 4 => "00000000"),
            217 => (0 => "11011001", 1 => "11011001", 2 => "11011001", 3 => "11011001", 4 => "00000000"),
            218 => (0 => "11011010", 1 => "11011010", 2 => "11011010", 3 => "11011010", 4 => "00000000"),
            219 => (0 => "11011011", 1 => "11011011", 2 => "11011011", 3 => "11011011", 4 => "00000000"),
            220 => (0 => "11011100", 1 => "11011100", 2 => "11011100", 3 => "11011100", 4 => "00000000"),
            221 => (0 => "11011101", 1 => "11011101", 2 => "11011101", 3 => "11011101", 4 => "00000000"),
            222 => (0 => "11011110", 1 => "11011110", 2 => "11011110", 3 => "11011110", 4 => "00000000"),
            223 => (0 => "11011111", 1 => "11011111", 2 => "11011111", 3 => "11011111", 4 => "00000000"),
            224 => (0 => "11100000", 1 => "11100000", 2 => "11100000", 3 => "11100000", 4 => "00000000"),
            225 => (0 => "11100001", 1 => "11100001", 2 => "11100001", 3 => "11100001", 4 => "00000000"),
            226 => (0 => "11100010", 1 => "11100010", 2 => "11100010", 3 => "11100010", 4 => "00000000"),
            227 => (0 => "11100011", 1 => "11100011", 2 => "11100011", 3 => "11100011", 4 => "00000000"),
            228 => (0 => "11100100", 1 => "11100100", 2 => "11100100", 3 => "11100100", 4 => "00000000"),
            229 => (0 => "11100101", 1 => "11100101", 2 => "11100101", 3 => "11100101", 4 => "00000000"),
            230 => (0 => "11100110", 1 => "11100110", 2 => "11100110", 3 => "11100110", 4 => "00000000"),
            231 => (0 => "11100111", 1 => "11100111", 2 => "11100111", 3 => "11100111", 4 => "00000000"),
            232 => (0 => "11101000", 1 => "11101000", 2 => "11101000", 3 => "11101000", 4 => "00000000"),
            233 => (0 => "11101001", 1 => "11101001", 2 => "11101001", 3 => "11101001", 4 => "00000000"),
            234 => (0 => "11101010", 1 => "11101010", 2 => "11101010", 3 => "11101010", 4 => "00000000"),
            235 => (0 => "11101011", 1 => "11101011", 2 => "11101011", 3 => "11101011", 4 => "00000000"),
            236 => (0 => "11101100", 1 => "11101100", 2 => "11101100", 3 => "11101100", 4 => "00000000"),
            237 => (0 => "11101101", 1 => "11101101", 2 => "11101101", 3 => "11101101", 4 => "00000000"),
            238 => (0 => "11101110", 1 => "11101110", 2 => "11101110", 3 => "11101110", 4 => "00000000"),
            239 => (0 => "11101111", 1 => "11101111", 2 => "11101111", 3 => "11101111", 4 => "00000000"),
            240 => (0 => "11110000", 1 => "11110000", 2 => "11110000", 3 => "11110000", 4 => "00000000"),
            241 => (0 => "11110001", 1 => "11110001", 2 => "11110001", 3 => "11110001", 4 => "00000000"),
            242 => (0 => "11110010", 1 => "11110010", 2 => "11110010", 3 => "11110010", 4 => "00000000"),
            243 => (0 => "11110011", 1 => "11110011", 2 => "11110011", 3 => "11110011", 4 => "00000000"),
            244 => (0 => "11110100", 1 => "11110100", 2 => "11110100", 3 => "11110100", 4 => "00000000"),
            245 => (0 => "11110101", 1 => "11110101", 2 => "11110101", 3 => "11110101", 4 => "00000000"),
            246 => (0 => "11110110", 1 => "11110110", 2 => "11110110", 3 => "11110110", 4 => "00000000"),
            247 => (0 => "11110111", 1 => "11110111", 2 => "11110111", 3 => "11110111", 4 => "00000000"),
            248 => (0 => "11111000", 1 => "11111000", 2 => "11111000", 3 => "11111000", 4 => "00000000"),
            249 => (0 => "11111001", 1 => "11111001", 2 => "11111001", 3 => "11111001", 4 => "00000000"),
            250 => (0 => "11111010", 1 => "11111010", 2 => "11111010", 3 => "11111010", 4 => "00000000"),
            251 => (0 => "11111011", 1 => "11111011", 2 => "11111011", 3 => "11111011", 4 => "00000000"),
            252 => (0 => "11111100", 1 => "11111100", 2 => "11111100", 3 => "11111100", 4 => "00000000"),
            253 => (0 => "11111101", 1 => "11111101", 2 => "11111101", 3 => "11111101", 4 => "00000000"),
            254 => (0 => "11111110", 1 => "11111110", 2 => "11111110", 3 => "11111110", 4 => "00000000"),
            255 => (0 => "11111111", 1 => "11111111", 2 => "11111111", 3 => "11111111", 4 => "00000000"),
            256 => (0 => "10000000", 1 => "00000000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            257 => (0 => "01000000", 1 => "00000000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            258 => (0 => "00100000", 1 => "00000000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            259 => (0 => "00010000", 1 => "00000000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            260 => (0 => "00001000", 1 => "00000000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            261 => (0 => "00000100", 1 => "00000000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            262 => (0 => "00000010", 1 => "00000000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            263 => (0 => "00000001", 1 => "00000000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            264 => (0 => "10000001", 1 => "00000001", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            265 => (0 => "01000001", 1 => "00000001", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            266 => (0 => "00100001", 1 => "00000001", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            267 => (0 => "00010001", 1 => "00000001", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            268 => (0 => "00001001", 1 => "00000001", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            269 => (0 => "00000101", 1 => "00000001", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            270 => (0 => "00000011", 1 => "00000001", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            271 => (0 => "00000000", 1 => "00000001", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            272 => (0 => "10000010", 1 => "00000010", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            273 => (0 => "01000010", 1 => "00000010", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            274 => (0 => "00100010", 1 => "00000010", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            275 => (0 => "00010010", 1 => "00000010", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            276 => (0 => "00001010", 1 => "00000010", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            277 => (0 => "00000110", 1 => "00000010", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            278 => (0 => "00000000", 1 => "00000010", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            279 => (0 => "00000011", 1 => "00000010", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            280 => (0 => "10000011", 1 => "00000011", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            281 => (0 => "01000011", 1 => "00000011", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            282 => (0 => "00100011", 1 => "00000011", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            283 => (0 => "00010011", 1 => "00000011", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            284 => (0 => "00001011", 1 => "00000011", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            285 => (0 => "00000111", 1 => "00000011", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            286 => (0 => "00000001", 1 => "00000011", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            287 => (0 => "00000010", 1 => "00000011", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            288 => (0 => "10000100", 1 => "00000100", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            289 => (0 => "01000100", 1 => "00000100", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            290 => (0 => "00100100", 1 => "00000100", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            291 => (0 => "00010100", 1 => "00000100", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            292 => (0 => "00001100", 1 => "00000100", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            293 => (0 => "00000000", 1 => "00000100", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            294 => (0 => "00000110", 1 => "00000100", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            295 => (0 => "00000101", 1 => "00000100", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            296 => (0 => "10000101", 1 => "00000101", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            297 => (0 => "01000101", 1 => "00000101", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            298 => (0 => "00100101", 1 => "00000101", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            299 => (0 => "00010101", 1 => "00000101", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            300 => (0 => "00001101", 1 => "00000101", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            301 => (0 => "00000001", 1 => "00000101", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            302 => (0 => "00000111", 1 => "00000101", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            303 => (0 => "00000100", 1 => "00000101", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            304 => (0 => "10000110", 1 => "00000110", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            305 => (0 => "01000110", 1 => "00000110", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            306 => (0 => "00100110", 1 => "00000110", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            307 => (0 => "00010110", 1 => "00000110", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            308 => (0 => "00001110", 1 => "00000110", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            309 => (0 => "00000010", 1 => "00000110", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            310 => (0 => "00000100", 1 => "00000110", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            311 => (0 => "00000111", 1 => "00000110", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            312 => (0 => "10000111", 1 => "00000111", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            313 => (0 => "01000111", 1 => "00000111", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            314 => (0 => "00100111", 1 => "00000111", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            315 => (0 => "00010111", 1 => "00000111", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            316 => (0 => "00001111", 1 => "00000111", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            317 => (0 => "00000011", 1 => "00000111", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            318 => (0 => "00000101", 1 => "00000111", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            319 => (0 => "00000110", 1 => "00000111", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            320 => (0 => "10001000", 1 => "00001000", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            321 => (0 => "01001000", 1 => "00001000", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            322 => (0 => "00101000", 1 => "00001000", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            323 => (0 => "00011000", 1 => "00001000", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            324 => (0 => "00000000", 1 => "00001000", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            325 => (0 => "00001100", 1 => "00001000", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            326 => (0 => "00001010", 1 => "00001000", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            327 => (0 => "00001001", 1 => "00001000", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            328 => (0 => "10001001", 1 => "00001001", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            329 => (0 => "01001001", 1 => "00001001", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            330 => (0 => "00101001", 1 => "00001001", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            331 => (0 => "00011001", 1 => "00001001", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            332 => (0 => "00000001", 1 => "00001001", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            333 => (0 => "00001101", 1 => "00001001", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            334 => (0 => "00001011", 1 => "00001001", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            335 => (0 => "00001000", 1 => "00001001", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            336 => (0 => "10001010", 1 => "00001010", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            337 => (0 => "01001010", 1 => "00001010", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            338 => (0 => "00101010", 1 => "00001010", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            339 => (0 => "00011010", 1 => "00001010", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            340 => (0 => "00000010", 1 => "00001010", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            341 => (0 => "00001110", 1 => "00001010", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            342 => (0 => "00001000", 1 => "00001010", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            343 => (0 => "00001011", 1 => "00001010", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            344 => (0 => "10001011", 1 => "00001011", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            345 => (0 => "01001011", 1 => "00001011", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            346 => (0 => "00101011", 1 => "00001011", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            347 => (0 => "00011011", 1 => "00001011", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            348 => (0 => "00000011", 1 => "00001011", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            349 => (0 => "00001111", 1 => "00001011", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            350 => (0 => "00001001", 1 => "00001011", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            351 => (0 => "00001010", 1 => "00001011", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            352 => (0 => "10001100", 1 => "00001100", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            353 => (0 => "01001100", 1 => "00001100", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            354 => (0 => "00101100", 1 => "00001100", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            355 => (0 => "00011100", 1 => "00001100", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            356 => (0 => "00000100", 1 => "00001100", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            357 => (0 => "00001000", 1 => "00001100", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            358 => (0 => "00001110", 1 => "00001100", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            359 => (0 => "00001101", 1 => "00001100", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            360 => (0 => "10001101", 1 => "00001101", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            361 => (0 => "01001101", 1 => "00001101", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            362 => (0 => "00101101", 1 => "00001101", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            363 => (0 => "00011101", 1 => "00001101", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            364 => (0 => "00000101", 1 => "00001101", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            365 => (0 => "00001001", 1 => "00001101", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            366 => (0 => "00001111", 1 => "00001101", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            367 => (0 => "00001100", 1 => "00001101", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            368 => (0 => "10001110", 1 => "00001110", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            369 => (0 => "01001110", 1 => "00001110", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            370 => (0 => "00101110", 1 => "00001110", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            371 => (0 => "00011110", 1 => "00001110", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            372 => (0 => "00000110", 1 => "00001110", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            373 => (0 => "00001010", 1 => "00001110", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            374 => (0 => "00001100", 1 => "00001110", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            375 => (0 => "00001111", 1 => "00001110", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            376 => (0 => "10001111", 1 => "00001111", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            377 => (0 => "01001111", 1 => "00001111", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            378 => (0 => "00101111", 1 => "00001111", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            379 => (0 => "00011111", 1 => "00001111", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            380 => (0 => "00000111", 1 => "00001111", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            381 => (0 => "00001011", 1 => "00001111", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            382 => (0 => "00001101", 1 => "00001111", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            383 => (0 => "00001110", 1 => "00001111", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            384 => (0 => "10010000", 1 => "00010000", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            385 => (0 => "01010000", 1 => "00010000", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            386 => (0 => "00110000", 1 => "00010000", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            387 => (0 => "00000000", 1 => "00010000", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            388 => (0 => "00011000", 1 => "00010000", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            389 => (0 => "00010100", 1 => "00010000", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            390 => (0 => "00010010", 1 => "00010000", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            391 => (0 => "00010001", 1 => "00010000", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            392 => (0 => "10010001", 1 => "00010001", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            393 => (0 => "01010001", 1 => "00010001", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            394 => (0 => "00110001", 1 => "00010001", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            395 => (0 => "00000001", 1 => "00010001", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            396 => (0 => "00011001", 1 => "00010001", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            397 => (0 => "00010101", 1 => "00010001", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            398 => (0 => "00010011", 1 => "00010001", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            399 => (0 => "00010000", 1 => "00010001", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            400 => (0 => "10010010", 1 => "00010010", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            401 => (0 => "01010010", 1 => "00010010", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            402 => (0 => "00110010", 1 => "00010010", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            403 => (0 => "00000010", 1 => "00010010", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            404 => (0 => "00011010", 1 => "00010010", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            405 => (0 => "00010110", 1 => "00010010", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            406 => (0 => "00010000", 1 => "00010010", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            407 => (0 => "00010011", 1 => "00010010", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            408 => (0 => "10010011", 1 => "00010011", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            409 => (0 => "01010011", 1 => "00010011", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            410 => (0 => "00110011", 1 => "00010011", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            411 => (0 => "00000011", 1 => "00010011", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            412 => (0 => "00011011", 1 => "00010011", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            413 => (0 => "00010111", 1 => "00010011", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            414 => (0 => "00010001", 1 => "00010011", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            415 => (0 => "00010010", 1 => "00010011", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            416 => (0 => "10010100", 1 => "00010100", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            417 => (0 => "01010100", 1 => "00010100", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            418 => (0 => "00110100", 1 => "00010100", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            419 => (0 => "00000100", 1 => "00010100", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            420 => (0 => "00011100", 1 => "00010100", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            421 => (0 => "00010000", 1 => "00010100", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            422 => (0 => "00010110", 1 => "00010100", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            423 => (0 => "00010101", 1 => "00010100", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            424 => (0 => "10010101", 1 => "00010101", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            425 => (0 => "01010101", 1 => "00010101", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            426 => (0 => "00110101", 1 => "00010101", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            427 => (0 => "00000101", 1 => "00010101", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            428 => (0 => "00011101", 1 => "00010101", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            429 => (0 => "00010001", 1 => "00010101", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            430 => (0 => "00010111", 1 => "00010101", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            431 => (0 => "00010100", 1 => "00010101", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            432 => (0 => "10010110", 1 => "00010110", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            433 => (0 => "01010110", 1 => "00010110", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            434 => (0 => "00110110", 1 => "00010110", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            435 => (0 => "00000110", 1 => "00010110", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            436 => (0 => "00011110", 1 => "00010110", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            437 => (0 => "00010010", 1 => "00010110", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            438 => (0 => "00010100", 1 => "00010110", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            439 => (0 => "00010111", 1 => "00010110", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            440 => (0 => "10010111", 1 => "00010111", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            441 => (0 => "01010111", 1 => "00010111", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            442 => (0 => "00110111", 1 => "00010111", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            443 => (0 => "00000111", 1 => "00010111", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            444 => (0 => "00011111", 1 => "00010111", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            445 => (0 => "00010011", 1 => "00010111", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            446 => (0 => "00010101", 1 => "00010111", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            447 => (0 => "00010110", 1 => "00010111", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            448 => (0 => "10011000", 1 => "00011000", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            449 => (0 => "01011000", 1 => "00011000", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            450 => (0 => "00111000", 1 => "00011000", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            451 => (0 => "00001000", 1 => "00011000", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            452 => (0 => "00010000", 1 => "00011000", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            453 => (0 => "00011100", 1 => "00011000", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            454 => (0 => "00011010", 1 => "00011000", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            455 => (0 => "00011001", 1 => "00011000", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            456 => (0 => "10011001", 1 => "00011001", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            457 => (0 => "01011001", 1 => "00011001", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            458 => (0 => "00111001", 1 => "00011001", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            459 => (0 => "00001001", 1 => "00011001", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            460 => (0 => "00010001", 1 => "00011001", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            461 => (0 => "00011101", 1 => "00011001", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            462 => (0 => "00011011", 1 => "00011001", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            463 => (0 => "00011000", 1 => "00011001", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            464 => (0 => "10011010", 1 => "00011010", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            465 => (0 => "01011010", 1 => "00011010", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            466 => (0 => "00111010", 1 => "00011010", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            467 => (0 => "00001010", 1 => "00011010", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            468 => (0 => "00010010", 1 => "00011010", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            469 => (0 => "00011110", 1 => "00011010", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            470 => (0 => "00011000", 1 => "00011010", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            471 => (0 => "00011011", 1 => "00011010", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            472 => (0 => "10011011", 1 => "00011011", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            473 => (0 => "01011011", 1 => "00011011", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            474 => (0 => "00111011", 1 => "00011011", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            475 => (0 => "00001011", 1 => "00011011", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            476 => (0 => "00010011", 1 => "00011011", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            477 => (0 => "00011111", 1 => "00011011", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            478 => (0 => "00011001", 1 => "00011011", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            479 => (0 => "00011010", 1 => "00011011", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            480 => (0 => "10011100", 1 => "00011100", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            481 => (0 => "01011100", 1 => "00011100", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            482 => (0 => "00111100", 1 => "00011100", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            483 => (0 => "00001100", 1 => "00011100", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            484 => (0 => "00010100", 1 => "00011100", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            485 => (0 => "00011000", 1 => "00011100", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            486 => (0 => "00011110", 1 => "00011100", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            487 => (0 => "00011101", 1 => "00011100", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            488 => (0 => "10011101", 1 => "00011101", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            489 => (0 => "01011101", 1 => "00011101", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            490 => (0 => "00111101", 1 => "00011101", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            491 => (0 => "00001101", 1 => "00011101", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            492 => (0 => "00010101", 1 => "00011101", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            493 => (0 => "00011001", 1 => "00011101", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            494 => (0 => "00011111", 1 => "00011101", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            495 => (0 => "00011100", 1 => "00011101", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            496 => (0 => "10011110", 1 => "00011110", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            497 => (0 => "01011110", 1 => "00011110", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            498 => (0 => "00111110", 1 => "00011110", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            499 => (0 => "00001110", 1 => "00011110", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            500 => (0 => "00010110", 1 => "00011110", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            501 => (0 => "00011010", 1 => "00011110", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            502 => (0 => "00011100", 1 => "00011110", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            503 => (0 => "00011111", 1 => "00011110", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            504 => (0 => "10011111", 1 => "00011111", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            505 => (0 => "01011111", 1 => "00011111", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            506 => (0 => "00111111", 1 => "00011111", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            507 => (0 => "00001111", 1 => "00011111", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            508 => (0 => "00010111", 1 => "00011111", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            509 => (0 => "00011011", 1 => "00011111", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            510 => (0 => "00011101", 1 => "00011111", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            511 => (0 => "00011110", 1 => "00011111", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            512 => (0 => "10100000", 1 => "00100000", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            513 => (0 => "01100000", 1 => "00100000", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            514 => (0 => "00000000", 1 => "00100000", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            515 => (0 => "00110000", 1 => "00100000", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            516 => (0 => "00101000", 1 => "00100000", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            517 => (0 => "00100100", 1 => "00100000", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            518 => (0 => "00100010", 1 => "00100000", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            519 => (0 => "00100001", 1 => "00100000", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            520 => (0 => "10100001", 1 => "00100001", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            521 => (0 => "01100001", 1 => "00100001", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            522 => (0 => "00000001", 1 => "00100001", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            523 => (0 => "00110001", 1 => "00100001", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            524 => (0 => "00101001", 1 => "00100001", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            525 => (0 => "00100101", 1 => "00100001", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            526 => (0 => "00100011", 1 => "00100001", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            527 => (0 => "00100000", 1 => "00100001", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            528 => (0 => "10100010", 1 => "00100010", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            529 => (0 => "01100010", 1 => "00100010", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            530 => (0 => "00000010", 1 => "00100010", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            531 => (0 => "00110010", 1 => "00100010", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            532 => (0 => "00101010", 1 => "00100010", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            533 => (0 => "00100110", 1 => "00100010", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            534 => (0 => "00100000", 1 => "00100010", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            535 => (0 => "00100011", 1 => "00100010", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            536 => (0 => "10100011", 1 => "00100011", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            537 => (0 => "01100011", 1 => "00100011", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            538 => (0 => "00000011", 1 => "00100011", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            539 => (0 => "00110011", 1 => "00100011", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            540 => (0 => "00101011", 1 => "00100011", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            541 => (0 => "00100111", 1 => "00100011", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            542 => (0 => "00100001", 1 => "00100011", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            543 => (0 => "00100010", 1 => "00100011", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            544 => (0 => "10100100", 1 => "00100100", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            545 => (0 => "01100100", 1 => "00100100", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            546 => (0 => "00000100", 1 => "00100100", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            547 => (0 => "00110100", 1 => "00100100", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            548 => (0 => "00101100", 1 => "00100100", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            549 => (0 => "00100000", 1 => "00100100", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            550 => (0 => "00100110", 1 => "00100100", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            551 => (0 => "00100101", 1 => "00100100", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            552 => (0 => "10100101", 1 => "00100101", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            553 => (0 => "01100101", 1 => "00100101", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            554 => (0 => "00000101", 1 => "00100101", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            555 => (0 => "00110101", 1 => "00100101", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            556 => (0 => "00101101", 1 => "00100101", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            557 => (0 => "00100001", 1 => "00100101", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            558 => (0 => "00100111", 1 => "00100101", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            559 => (0 => "00100100", 1 => "00100101", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            560 => (0 => "10100110", 1 => "00100110", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            561 => (0 => "01100110", 1 => "00100110", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            562 => (0 => "00000110", 1 => "00100110", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            563 => (0 => "00110110", 1 => "00100110", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            564 => (0 => "00101110", 1 => "00100110", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            565 => (0 => "00100010", 1 => "00100110", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            566 => (0 => "00100100", 1 => "00100110", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            567 => (0 => "00100111", 1 => "00100110", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            568 => (0 => "10100111", 1 => "00100111", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            569 => (0 => "01100111", 1 => "00100111", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            570 => (0 => "00000111", 1 => "00100111", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            571 => (0 => "00110111", 1 => "00100111", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            572 => (0 => "00101111", 1 => "00100111", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            573 => (0 => "00100011", 1 => "00100111", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            574 => (0 => "00100101", 1 => "00100111", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            575 => (0 => "00100110", 1 => "00100111", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            576 => (0 => "10101000", 1 => "00101000", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            577 => (0 => "01101000", 1 => "00101000", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            578 => (0 => "00001000", 1 => "00101000", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            579 => (0 => "00111000", 1 => "00101000", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            580 => (0 => "00100000", 1 => "00101000", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            581 => (0 => "00101100", 1 => "00101000", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            582 => (0 => "00101010", 1 => "00101000", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            583 => (0 => "00101001", 1 => "00101000", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            584 => (0 => "10101001", 1 => "00101001", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            585 => (0 => "01101001", 1 => "00101001", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            586 => (0 => "00001001", 1 => "00101001", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            587 => (0 => "00111001", 1 => "00101001", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            588 => (0 => "00100001", 1 => "00101001", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            589 => (0 => "00101101", 1 => "00101001", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            590 => (0 => "00101011", 1 => "00101001", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            591 => (0 => "00101000", 1 => "00101001", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            592 => (0 => "10101010", 1 => "00101010", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            593 => (0 => "01101010", 1 => "00101010", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            594 => (0 => "00001010", 1 => "00101010", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            595 => (0 => "00111010", 1 => "00101010", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            596 => (0 => "00100010", 1 => "00101010", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            597 => (0 => "00101110", 1 => "00101010", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            598 => (0 => "00101000", 1 => "00101010", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            599 => (0 => "00101011", 1 => "00101010", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            600 => (0 => "10101011", 1 => "00101011", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            601 => (0 => "01101011", 1 => "00101011", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            602 => (0 => "00001011", 1 => "00101011", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            603 => (0 => "00111011", 1 => "00101011", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            604 => (0 => "00100011", 1 => "00101011", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            605 => (0 => "00101111", 1 => "00101011", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            606 => (0 => "00101001", 1 => "00101011", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            607 => (0 => "00101010", 1 => "00101011", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            608 => (0 => "10101100", 1 => "00101100", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            609 => (0 => "01101100", 1 => "00101100", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            610 => (0 => "00001100", 1 => "00101100", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            611 => (0 => "00111100", 1 => "00101100", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            612 => (0 => "00100100", 1 => "00101100", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            613 => (0 => "00101000", 1 => "00101100", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            614 => (0 => "00101110", 1 => "00101100", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            615 => (0 => "00101101", 1 => "00101100", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            616 => (0 => "10101101", 1 => "00101101", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            617 => (0 => "01101101", 1 => "00101101", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            618 => (0 => "00001101", 1 => "00101101", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            619 => (0 => "00111101", 1 => "00101101", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            620 => (0 => "00100101", 1 => "00101101", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            621 => (0 => "00101001", 1 => "00101101", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            622 => (0 => "00101111", 1 => "00101101", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            623 => (0 => "00101100", 1 => "00101101", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            624 => (0 => "10101110", 1 => "00101110", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            625 => (0 => "01101110", 1 => "00101110", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            626 => (0 => "00001110", 1 => "00101110", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            627 => (0 => "00111110", 1 => "00101110", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            628 => (0 => "00100110", 1 => "00101110", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            629 => (0 => "00101010", 1 => "00101110", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            630 => (0 => "00101100", 1 => "00101110", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            631 => (0 => "00101111", 1 => "00101110", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            632 => (0 => "10101111", 1 => "00101111", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            633 => (0 => "01101111", 1 => "00101111", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            634 => (0 => "00001111", 1 => "00101111", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            635 => (0 => "00111111", 1 => "00101111", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            636 => (0 => "00100111", 1 => "00101111", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            637 => (0 => "00101011", 1 => "00101111", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            638 => (0 => "00101101", 1 => "00101111", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            639 => (0 => "00101110", 1 => "00101111", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            640 => (0 => "10110000", 1 => "00110000", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            641 => (0 => "01110000", 1 => "00110000", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            642 => (0 => "00010000", 1 => "00110000", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            643 => (0 => "00100000", 1 => "00110000", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            644 => (0 => "00111000", 1 => "00110000", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            645 => (0 => "00110100", 1 => "00110000", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            646 => (0 => "00110010", 1 => "00110000", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            647 => (0 => "00110001", 1 => "00110000", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            648 => (0 => "10110001", 1 => "00110001", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            649 => (0 => "01110001", 1 => "00110001", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            650 => (0 => "00010001", 1 => "00110001", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            651 => (0 => "00100001", 1 => "00110001", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            652 => (0 => "00111001", 1 => "00110001", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            653 => (0 => "00110101", 1 => "00110001", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            654 => (0 => "00110011", 1 => "00110001", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            655 => (0 => "00110000", 1 => "00110001", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            656 => (0 => "10110010", 1 => "00110010", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            657 => (0 => "01110010", 1 => "00110010", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            658 => (0 => "00010010", 1 => "00110010", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            659 => (0 => "00100010", 1 => "00110010", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            660 => (0 => "00111010", 1 => "00110010", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            661 => (0 => "00110110", 1 => "00110010", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            662 => (0 => "00110000", 1 => "00110010", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            663 => (0 => "00110011", 1 => "00110010", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            664 => (0 => "10110011", 1 => "00110011", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            665 => (0 => "01110011", 1 => "00110011", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            666 => (0 => "00010011", 1 => "00110011", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            667 => (0 => "00100011", 1 => "00110011", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            668 => (0 => "00111011", 1 => "00110011", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            669 => (0 => "00110111", 1 => "00110011", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            670 => (0 => "00110001", 1 => "00110011", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            671 => (0 => "00110010", 1 => "00110011", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            672 => (0 => "10110100", 1 => "00110100", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            673 => (0 => "01110100", 1 => "00110100", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            674 => (0 => "00010100", 1 => "00110100", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            675 => (0 => "00100100", 1 => "00110100", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            676 => (0 => "00111100", 1 => "00110100", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            677 => (0 => "00110000", 1 => "00110100", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            678 => (0 => "00110110", 1 => "00110100", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            679 => (0 => "00110101", 1 => "00110100", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            680 => (0 => "10110101", 1 => "00110101", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            681 => (0 => "01110101", 1 => "00110101", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            682 => (0 => "00010101", 1 => "00110101", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            683 => (0 => "00100101", 1 => "00110101", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            684 => (0 => "00111101", 1 => "00110101", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            685 => (0 => "00110001", 1 => "00110101", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            686 => (0 => "00110111", 1 => "00110101", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            687 => (0 => "00110100", 1 => "00110101", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            688 => (0 => "10110110", 1 => "00110110", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            689 => (0 => "01110110", 1 => "00110110", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            690 => (0 => "00010110", 1 => "00110110", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            691 => (0 => "00100110", 1 => "00110110", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            692 => (0 => "00111110", 1 => "00110110", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            693 => (0 => "00110010", 1 => "00110110", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            694 => (0 => "00110100", 1 => "00110110", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            695 => (0 => "00110111", 1 => "00110110", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            696 => (0 => "10110111", 1 => "00110111", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            697 => (0 => "01110111", 1 => "00110111", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            698 => (0 => "00010111", 1 => "00110111", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            699 => (0 => "00100111", 1 => "00110111", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            700 => (0 => "00111111", 1 => "00110111", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            701 => (0 => "00110011", 1 => "00110111", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            702 => (0 => "00110101", 1 => "00110111", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            703 => (0 => "00110110", 1 => "00110111", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            704 => (0 => "10111000", 1 => "00111000", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            705 => (0 => "01111000", 1 => "00111000", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            706 => (0 => "00011000", 1 => "00111000", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            707 => (0 => "00101000", 1 => "00111000", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            708 => (0 => "00110000", 1 => "00111000", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            709 => (0 => "00111100", 1 => "00111000", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            710 => (0 => "00111010", 1 => "00111000", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            711 => (0 => "00111001", 1 => "00111000", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            712 => (0 => "10111001", 1 => "00111001", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            713 => (0 => "01111001", 1 => "00111001", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            714 => (0 => "00011001", 1 => "00111001", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            715 => (0 => "00101001", 1 => "00111001", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            716 => (0 => "00110001", 1 => "00111001", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            717 => (0 => "00111101", 1 => "00111001", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            718 => (0 => "00111011", 1 => "00111001", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            719 => (0 => "00111000", 1 => "00111001", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            720 => (0 => "10111010", 1 => "00111010", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            721 => (0 => "01111010", 1 => "00111010", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            722 => (0 => "00011010", 1 => "00111010", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            723 => (0 => "00101010", 1 => "00111010", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            724 => (0 => "00110010", 1 => "00111010", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            725 => (0 => "00111110", 1 => "00111010", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            726 => (0 => "00111000", 1 => "00111010", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            727 => (0 => "00111011", 1 => "00111010", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            728 => (0 => "10111011", 1 => "00111011", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            729 => (0 => "01111011", 1 => "00111011", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            730 => (0 => "00011011", 1 => "00111011", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            731 => (0 => "00101011", 1 => "00111011", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            732 => (0 => "00110011", 1 => "00111011", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            733 => (0 => "00111111", 1 => "00111011", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            734 => (0 => "00111001", 1 => "00111011", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            735 => (0 => "00111010", 1 => "00111011", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            736 => (0 => "10111100", 1 => "00111100", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            737 => (0 => "01111100", 1 => "00111100", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            738 => (0 => "00011100", 1 => "00111100", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            739 => (0 => "00101100", 1 => "00111100", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            740 => (0 => "00110100", 1 => "00111100", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            741 => (0 => "00111000", 1 => "00111100", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            742 => (0 => "00111110", 1 => "00111100", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            743 => (0 => "00111101", 1 => "00111100", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            744 => (0 => "10111101", 1 => "00111101", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            745 => (0 => "01111101", 1 => "00111101", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            746 => (0 => "00011101", 1 => "00111101", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            747 => (0 => "00101101", 1 => "00111101", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            748 => (0 => "00110101", 1 => "00111101", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            749 => (0 => "00111001", 1 => "00111101", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            750 => (0 => "00111111", 1 => "00111101", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            751 => (0 => "00111100", 1 => "00111101", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            752 => (0 => "10111110", 1 => "00111110", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            753 => (0 => "01111110", 1 => "00111110", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            754 => (0 => "00011110", 1 => "00111110", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            755 => (0 => "00101110", 1 => "00111110", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            756 => (0 => "00110110", 1 => "00111110", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            757 => (0 => "00111010", 1 => "00111110", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            758 => (0 => "00111100", 1 => "00111110", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            759 => (0 => "00111111", 1 => "00111110", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            760 => (0 => "10111111", 1 => "00111111", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            761 => (0 => "01111111", 1 => "00111111", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            762 => (0 => "00011111", 1 => "00111111", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            763 => (0 => "00101111", 1 => "00111111", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            764 => (0 => "00110111", 1 => "00111111", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            765 => (0 => "00111011", 1 => "00111111", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            766 => (0 => "00111101", 1 => "00111111", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            767 => (0 => "00111110", 1 => "00111111", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            768 => (0 => "11000000", 1 => "01000000", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            769 => (0 => "00000000", 1 => "01000000", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            770 => (0 => "01100000", 1 => "01000000", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            771 => (0 => "01010000", 1 => "01000000", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            772 => (0 => "01001000", 1 => "01000000", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            773 => (0 => "01000100", 1 => "01000000", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            774 => (0 => "01000010", 1 => "01000000", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            775 => (0 => "01000001", 1 => "01000000", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            776 => (0 => "11000001", 1 => "01000001", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            777 => (0 => "00000001", 1 => "01000001", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            778 => (0 => "01100001", 1 => "01000001", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            779 => (0 => "01010001", 1 => "01000001", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            780 => (0 => "01001001", 1 => "01000001", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            781 => (0 => "01000101", 1 => "01000001", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            782 => (0 => "01000011", 1 => "01000001", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            783 => (0 => "01000000", 1 => "01000001", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            784 => (0 => "11000010", 1 => "01000010", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            785 => (0 => "00000010", 1 => "01000010", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            786 => (0 => "01100010", 1 => "01000010", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            787 => (0 => "01010010", 1 => "01000010", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            788 => (0 => "01001010", 1 => "01000010", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            789 => (0 => "01000110", 1 => "01000010", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            790 => (0 => "01000000", 1 => "01000010", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            791 => (0 => "01000011", 1 => "01000010", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            792 => (0 => "11000011", 1 => "01000011", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            793 => (0 => "00000011", 1 => "01000011", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            794 => (0 => "01100011", 1 => "01000011", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            795 => (0 => "01010011", 1 => "01000011", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            796 => (0 => "01001011", 1 => "01000011", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            797 => (0 => "01000111", 1 => "01000011", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            798 => (0 => "01000001", 1 => "01000011", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            799 => (0 => "01000010", 1 => "01000011", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            800 => (0 => "11000100", 1 => "01000100", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            801 => (0 => "00000100", 1 => "01000100", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            802 => (0 => "01100100", 1 => "01000100", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            803 => (0 => "01010100", 1 => "01000100", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            804 => (0 => "01001100", 1 => "01000100", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            805 => (0 => "01000000", 1 => "01000100", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            806 => (0 => "01000110", 1 => "01000100", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            807 => (0 => "01000101", 1 => "01000100", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            808 => (0 => "11000101", 1 => "01000101", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            809 => (0 => "00000101", 1 => "01000101", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            810 => (0 => "01100101", 1 => "01000101", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            811 => (0 => "01010101", 1 => "01000101", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            812 => (0 => "01001101", 1 => "01000101", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            813 => (0 => "01000001", 1 => "01000101", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            814 => (0 => "01000111", 1 => "01000101", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            815 => (0 => "01000100", 1 => "01000101", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            816 => (0 => "11000110", 1 => "01000110", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            817 => (0 => "00000110", 1 => "01000110", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            818 => (0 => "01100110", 1 => "01000110", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            819 => (0 => "01010110", 1 => "01000110", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            820 => (0 => "01001110", 1 => "01000110", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            821 => (0 => "01000010", 1 => "01000110", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            822 => (0 => "01000100", 1 => "01000110", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            823 => (0 => "01000111", 1 => "01000110", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            824 => (0 => "11000111", 1 => "01000111", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            825 => (0 => "00000111", 1 => "01000111", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            826 => (0 => "01100111", 1 => "01000111", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            827 => (0 => "01010111", 1 => "01000111", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            828 => (0 => "01001111", 1 => "01000111", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            829 => (0 => "01000011", 1 => "01000111", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            830 => (0 => "01000101", 1 => "01000111", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            831 => (0 => "01000110", 1 => "01000111", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            832 => (0 => "11001000", 1 => "01001000", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            833 => (0 => "00001000", 1 => "01001000", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            834 => (0 => "01101000", 1 => "01001000", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            835 => (0 => "01011000", 1 => "01001000", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            836 => (0 => "01000000", 1 => "01001000", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            837 => (0 => "01001100", 1 => "01001000", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            838 => (0 => "01001010", 1 => "01001000", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            839 => (0 => "01001001", 1 => "01001000", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            840 => (0 => "11001001", 1 => "01001001", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            841 => (0 => "00001001", 1 => "01001001", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            842 => (0 => "01101001", 1 => "01001001", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            843 => (0 => "01011001", 1 => "01001001", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            844 => (0 => "01000001", 1 => "01001001", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            845 => (0 => "01001101", 1 => "01001001", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            846 => (0 => "01001011", 1 => "01001001", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            847 => (0 => "01001000", 1 => "01001001", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            848 => (0 => "11001010", 1 => "01001010", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            849 => (0 => "00001010", 1 => "01001010", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            850 => (0 => "01101010", 1 => "01001010", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            851 => (0 => "01011010", 1 => "01001010", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            852 => (0 => "01000010", 1 => "01001010", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            853 => (0 => "01001110", 1 => "01001010", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            854 => (0 => "01001000", 1 => "01001010", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            855 => (0 => "01001011", 1 => "01001010", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            856 => (0 => "11001011", 1 => "01001011", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            857 => (0 => "00001011", 1 => "01001011", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            858 => (0 => "01101011", 1 => "01001011", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            859 => (0 => "01011011", 1 => "01001011", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            860 => (0 => "01000011", 1 => "01001011", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            861 => (0 => "01001111", 1 => "01001011", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            862 => (0 => "01001001", 1 => "01001011", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            863 => (0 => "01001010", 1 => "01001011", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            864 => (0 => "11001100", 1 => "01001100", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            865 => (0 => "00001100", 1 => "01001100", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            866 => (0 => "01101100", 1 => "01001100", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            867 => (0 => "01011100", 1 => "01001100", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            868 => (0 => "01000100", 1 => "01001100", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            869 => (0 => "01001000", 1 => "01001100", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            870 => (0 => "01001110", 1 => "01001100", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            871 => (0 => "01001101", 1 => "01001100", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            872 => (0 => "11001101", 1 => "01001101", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            873 => (0 => "00001101", 1 => "01001101", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            874 => (0 => "01101101", 1 => "01001101", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            875 => (0 => "01011101", 1 => "01001101", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            876 => (0 => "01000101", 1 => "01001101", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            877 => (0 => "01001001", 1 => "01001101", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            878 => (0 => "01001111", 1 => "01001101", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            879 => (0 => "01001100", 1 => "01001101", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            880 => (0 => "11001110", 1 => "01001110", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            881 => (0 => "00001110", 1 => "01001110", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            882 => (0 => "01101110", 1 => "01001110", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            883 => (0 => "01011110", 1 => "01001110", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            884 => (0 => "01000110", 1 => "01001110", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            885 => (0 => "01001010", 1 => "01001110", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            886 => (0 => "01001100", 1 => "01001110", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            887 => (0 => "01001111", 1 => "01001110", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            888 => (0 => "11001111", 1 => "01001111", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            889 => (0 => "00001111", 1 => "01001111", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            890 => (0 => "01101111", 1 => "01001111", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            891 => (0 => "01011111", 1 => "01001111", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            892 => (0 => "01000111", 1 => "01001111", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            893 => (0 => "01001011", 1 => "01001111", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            894 => (0 => "01001101", 1 => "01001111", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            895 => (0 => "01001110", 1 => "01001111", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            896 => (0 => "11010000", 1 => "01010000", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            897 => (0 => "00010000", 1 => "01010000", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            898 => (0 => "01110000", 1 => "01010000", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            899 => (0 => "01000000", 1 => "01010000", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            900 => (0 => "01011000", 1 => "01010000", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            901 => (0 => "01010100", 1 => "01010000", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            902 => (0 => "01010010", 1 => "01010000", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            903 => (0 => "01010001", 1 => "01010000", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            904 => (0 => "11010001", 1 => "01010001", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            905 => (0 => "00010001", 1 => "01010001", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            906 => (0 => "01110001", 1 => "01010001", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            907 => (0 => "01000001", 1 => "01010001", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            908 => (0 => "01011001", 1 => "01010001", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            909 => (0 => "01010101", 1 => "01010001", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            910 => (0 => "01010011", 1 => "01010001", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            911 => (0 => "01010000", 1 => "01010001", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            912 => (0 => "11010010", 1 => "01010010", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            913 => (0 => "00010010", 1 => "01010010", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            914 => (0 => "01110010", 1 => "01010010", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            915 => (0 => "01000010", 1 => "01010010", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            916 => (0 => "01011010", 1 => "01010010", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            917 => (0 => "01010110", 1 => "01010010", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            918 => (0 => "01010000", 1 => "01010010", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            919 => (0 => "01010011", 1 => "01010010", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            920 => (0 => "11010011", 1 => "01010011", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            921 => (0 => "00010011", 1 => "01010011", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            922 => (0 => "01110011", 1 => "01010011", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            923 => (0 => "01000011", 1 => "01010011", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            924 => (0 => "01011011", 1 => "01010011", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            925 => (0 => "01010111", 1 => "01010011", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            926 => (0 => "01010001", 1 => "01010011", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            927 => (0 => "01010010", 1 => "01010011", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            928 => (0 => "11010100", 1 => "01010100", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            929 => (0 => "00010100", 1 => "01010100", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            930 => (0 => "01110100", 1 => "01010100", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            931 => (0 => "01000100", 1 => "01010100", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            932 => (0 => "01011100", 1 => "01010100", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            933 => (0 => "01010000", 1 => "01010100", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            934 => (0 => "01010110", 1 => "01010100", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            935 => (0 => "01010101", 1 => "01010100", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            936 => (0 => "11010101", 1 => "01010101", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            937 => (0 => "00010101", 1 => "01010101", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            938 => (0 => "01110101", 1 => "01010101", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            939 => (0 => "01000101", 1 => "01010101", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            940 => (0 => "01011101", 1 => "01010101", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            941 => (0 => "01010001", 1 => "01010101", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            942 => (0 => "01010111", 1 => "01010101", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            943 => (0 => "01010100", 1 => "01010101", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            944 => (0 => "11010110", 1 => "01010110", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            945 => (0 => "00010110", 1 => "01010110", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            946 => (0 => "01110110", 1 => "01010110", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            947 => (0 => "01000110", 1 => "01010110", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            948 => (0 => "01011110", 1 => "01010110", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            949 => (0 => "01010010", 1 => "01010110", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            950 => (0 => "01010100", 1 => "01010110", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            951 => (0 => "01010111", 1 => "01010110", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            952 => (0 => "11010111", 1 => "01010111", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            953 => (0 => "00010111", 1 => "01010111", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            954 => (0 => "01110111", 1 => "01010111", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            955 => (0 => "01000111", 1 => "01010111", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            956 => (0 => "01011111", 1 => "01010111", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            957 => (0 => "01010011", 1 => "01010111", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            958 => (0 => "01010101", 1 => "01010111", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            959 => (0 => "01010110", 1 => "01010111", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            960 => (0 => "11011000", 1 => "01011000", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            961 => (0 => "00011000", 1 => "01011000", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            962 => (0 => "01111000", 1 => "01011000", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            963 => (0 => "01001000", 1 => "01011000", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            964 => (0 => "01010000", 1 => "01011000", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            965 => (0 => "01011100", 1 => "01011000", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            966 => (0 => "01011010", 1 => "01011000", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            967 => (0 => "01011001", 1 => "01011000", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            968 => (0 => "11011001", 1 => "01011001", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            969 => (0 => "00011001", 1 => "01011001", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            970 => (0 => "01111001", 1 => "01011001", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            971 => (0 => "01001001", 1 => "01011001", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            972 => (0 => "01010001", 1 => "01011001", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            973 => (0 => "01011101", 1 => "01011001", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            974 => (0 => "01011011", 1 => "01011001", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            975 => (0 => "01011000", 1 => "01011001", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            976 => (0 => "11011010", 1 => "01011010", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            977 => (0 => "00011010", 1 => "01011010", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            978 => (0 => "01111010", 1 => "01011010", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            979 => (0 => "01001010", 1 => "01011010", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            980 => (0 => "01010010", 1 => "01011010", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            981 => (0 => "01011110", 1 => "01011010", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            982 => (0 => "01011000", 1 => "01011010", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            983 => (0 => "01011011", 1 => "01011010", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            984 => (0 => "11011011", 1 => "01011011", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            985 => (0 => "00011011", 1 => "01011011", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            986 => (0 => "01111011", 1 => "01011011", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            987 => (0 => "01001011", 1 => "01011011", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            988 => (0 => "01010011", 1 => "01011011", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            989 => (0 => "01011111", 1 => "01011011", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            990 => (0 => "01011001", 1 => "01011011", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            991 => (0 => "01011010", 1 => "01011011", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            992 => (0 => "11011100", 1 => "01011100", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            993 => (0 => "00011100", 1 => "01011100", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            994 => (0 => "01111100", 1 => "01011100", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            995 => (0 => "01001100", 1 => "01011100", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            996 => (0 => "01010100", 1 => "01011100", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            997 => (0 => "01011000", 1 => "01011100", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            998 => (0 => "01011110", 1 => "01011100", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            999 => (0 => "01011101", 1 => "01011100", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            1000 => (0 => "11011101", 1 => "01011101", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            1001 => (0 => "00011101", 1 => "01011101", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            1002 => (0 => "01111101", 1 => "01011101", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            1003 => (0 => "01001101", 1 => "01011101", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            1004 => (0 => "01010101", 1 => "01011101", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            1005 => (0 => "01011001", 1 => "01011101", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            1006 => (0 => "01011111", 1 => "01011101", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            1007 => (0 => "01011100", 1 => "01011101", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            1008 => (0 => "11011110", 1 => "01011110", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            1009 => (0 => "00011110", 1 => "01011110", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            1010 => (0 => "01111110", 1 => "01011110", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            1011 => (0 => "01001110", 1 => "01011110", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            1012 => (0 => "01010110", 1 => "01011110", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            1013 => (0 => "01011010", 1 => "01011110", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            1014 => (0 => "01011100", 1 => "01011110", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            1015 => (0 => "01011111", 1 => "01011110", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            1016 => (0 => "11011111", 1 => "01011111", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            1017 => (0 => "00011111", 1 => "01011111", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            1018 => (0 => "01111111", 1 => "01011111", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            1019 => (0 => "01001111", 1 => "01011111", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            1020 => (0 => "01010111", 1 => "01011111", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            1021 => (0 => "01011011", 1 => "01011111", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            1022 => (0 => "01011101", 1 => "01011111", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            1023 => (0 => "01011110", 1 => "01011111", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            1024 => (0 => "11100000", 1 => "01100000", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            1025 => (0 => "00100000", 1 => "01100000", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            1026 => (0 => "01000000", 1 => "01100000", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            1027 => (0 => "01110000", 1 => "01100000", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            1028 => (0 => "01101000", 1 => "01100000", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            1029 => (0 => "01100100", 1 => "01100000", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            1030 => (0 => "01100010", 1 => "01100000", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            1031 => (0 => "01100001", 1 => "01100000", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            1032 => (0 => "11100001", 1 => "01100001", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            1033 => (0 => "00100001", 1 => "01100001", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            1034 => (0 => "01000001", 1 => "01100001", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            1035 => (0 => "01110001", 1 => "01100001", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            1036 => (0 => "01101001", 1 => "01100001", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            1037 => (0 => "01100101", 1 => "01100001", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            1038 => (0 => "01100011", 1 => "01100001", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            1039 => (0 => "01100000", 1 => "01100001", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            1040 => (0 => "11100010", 1 => "01100010", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            1041 => (0 => "00100010", 1 => "01100010", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            1042 => (0 => "01000010", 1 => "01100010", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            1043 => (0 => "01110010", 1 => "01100010", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            1044 => (0 => "01101010", 1 => "01100010", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            1045 => (0 => "01100110", 1 => "01100010", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            1046 => (0 => "01100000", 1 => "01100010", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            1047 => (0 => "01100011", 1 => "01100010", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            1048 => (0 => "11100011", 1 => "01100011", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            1049 => (0 => "00100011", 1 => "01100011", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            1050 => (0 => "01000011", 1 => "01100011", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            1051 => (0 => "01110011", 1 => "01100011", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            1052 => (0 => "01101011", 1 => "01100011", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            1053 => (0 => "01100111", 1 => "01100011", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            1054 => (0 => "01100001", 1 => "01100011", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            1055 => (0 => "01100010", 1 => "01100011", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            1056 => (0 => "11100100", 1 => "01100100", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            1057 => (0 => "00100100", 1 => "01100100", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            1058 => (0 => "01000100", 1 => "01100100", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            1059 => (0 => "01110100", 1 => "01100100", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            1060 => (0 => "01101100", 1 => "01100100", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            1061 => (0 => "01100000", 1 => "01100100", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            1062 => (0 => "01100110", 1 => "01100100", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            1063 => (0 => "01100101", 1 => "01100100", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            1064 => (0 => "11100101", 1 => "01100101", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            1065 => (0 => "00100101", 1 => "01100101", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            1066 => (0 => "01000101", 1 => "01100101", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            1067 => (0 => "01110101", 1 => "01100101", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            1068 => (0 => "01101101", 1 => "01100101", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            1069 => (0 => "01100001", 1 => "01100101", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            1070 => (0 => "01100111", 1 => "01100101", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            1071 => (0 => "01100100", 1 => "01100101", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            1072 => (0 => "11100110", 1 => "01100110", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            1073 => (0 => "00100110", 1 => "01100110", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            1074 => (0 => "01000110", 1 => "01100110", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            1075 => (0 => "01110110", 1 => "01100110", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            1076 => (0 => "01101110", 1 => "01100110", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            1077 => (0 => "01100010", 1 => "01100110", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            1078 => (0 => "01100100", 1 => "01100110", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            1079 => (0 => "01100111", 1 => "01100110", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            1080 => (0 => "11100111", 1 => "01100111", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            1081 => (0 => "00100111", 1 => "01100111", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            1082 => (0 => "01000111", 1 => "01100111", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            1083 => (0 => "01110111", 1 => "01100111", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            1084 => (0 => "01101111", 1 => "01100111", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            1085 => (0 => "01100011", 1 => "01100111", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            1086 => (0 => "01100101", 1 => "01100111", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            1087 => (0 => "01100110", 1 => "01100111", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            1088 => (0 => "11101000", 1 => "01101000", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            1089 => (0 => "00101000", 1 => "01101000", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            1090 => (0 => "01001000", 1 => "01101000", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            1091 => (0 => "01111000", 1 => "01101000", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            1092 => (0 => "01100000", 1 => "01101000", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            1093 => (0 => "01101100", 1 => "01101000", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            1094 => (0 => "01101010", 1 => "01101000", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            1095 => (0 => "01101001", 1 => "01101000", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            1096 => (0 => "11101001", 1 => "01101001", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            1097 => (0 => "00101001", 1 => "01101001", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            1098 => (0 => "01001001", 1 => "01101001", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            1099 => (0 => "01111001", 1 => "01101001", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            1100 => (0 => "01100001", 1 => "01101001", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            1101 => (0 => "01101101", 1 => "01101001", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            1102 => (0 => "01101011", 1 => "01101001", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            1103 => (0 => "01101000", 1 => "01101001", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            1104 => (0 => "11101010", 1 => "01101010", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            1105 => (0 => "00101010", 1 => "01101010", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            1106 => (0 => "01001010", 1 => "01101010", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            1107 => (0 => "01111010", 1 => "01101010", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            1108 => (0 => "01100010", 1 => "01101010", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            1109 => (0 => "01101110", 1 => "01101010", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            1110 => (0 => "01101000", 1 => "01101010", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            1111 => (0 => "01101011", 1 => "01101010", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            1112 => (0 => "11101011", 1 => "01101011", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            1113 => (0 => "00101011", 1 => "01101011", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            1114 => (0 => "01001011", 1 => "01101011", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            1115 => (0 => "01111011", 1 => "01101011", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            1116 => (0 => "01100011", 1 => "01101011", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            1117 => (0 => "01101111", 1 => "01101011", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            1118 => (0 => "01101001", 1 => "01101011", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            1119 => (0 => "01101010", 1 => "01101011", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            1120 => (0 => "11101100", 1 => "01101100", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            1121 => (0 => "00101100", 1 => "01101100", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            1122 => (0 => "01001100", 1 => "01101100", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            1123 => (0 => "01111100", 1 => "01101100", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            1124 => (0 => "01100100", 1 => "01101100", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            1125 => (0 => "01101000", 1 => "01101100", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            1126 => (0 => "01101110", 1 => "01101100", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            1127 => (0 => "01101101", 1 => "01101100", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            1128 => (0 => "11101101", 1 => "01101101", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            1129 => (0 => "00101101", 1 => "01101101", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            1130 => (0 => "01001101", 1 => "01101101", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            1131 => (0 => "01111101", 1 => "01101101", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            1132 => (0 => "01100101", 1 => "01101101", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            1133 => (0 => "01101001", 1 => "01101101", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            1134 => (0 => "01101111", 1 => "01101101", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            1135 => (0 => "01101100", 1 => "01101101", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            1136 => (0 => "11101110", 1 => "01101110", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            1137 => (0 => "00101110", 1 => "01101110", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            1138 => (0 => "01001110", 1 => "01101110", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            1139 => (0 => "01111110", 1 => "01101110", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            1140 => (0 => "01100110", 1 => "01101110", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            1141 => (0 => "01101010", 1 => "01101110", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            1142 => (0 => "01101100", 1 => "01101110", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            1143 => (0 => "01101111", 1 => "01101110", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            1144 => (0 => "11101111", 1 => "01101111", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            1145 => (0 => "00101111", 1 => "01101111", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            1146 => (0 => "01001111", 1 => "01101111", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            1147 => (0 => "01111111", 1 => "01101111", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            1148 => (0 => "01100111", 1 => "01101111", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            1149 => (0 => "01101011", 1 => "01101111", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            1150 => (0 => "01101101", 1 => "01101111", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            1151 => (0 => "01101110", 1 => "01101111", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            1152 => (0 => "11110000", 1 => "01110000", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            1153 => (0 => "00110000", 1 => "01110000", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            1154 => (0 => "01010000", 1 => "01110000", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            1155 => (0 => "01100000", 1 => "01110000", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            1156 => (0 => "01111000", 1 => "01110000", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            1157 => (0 => "01110100", 1 => "01110000", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            1158 => (0 => "01110010", 1 => "01110000", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            1159 => (0 => "01110001", 1 => "01110000", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            1160 => (0 => "11110001", 1 => "01110001", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            1161 => (0 => "00110001", 1 => "01110001", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            1162 => (0 => "01010001", 1 => "01110001", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            1163 => (0 => "01100001", 1 => "01110001", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            1164 => (0 => "01111001", 1 => "01110001", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            1165 => (0 => "01110101", 1 => "01110001", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            1166 => (0 => "01110011", 1 => "01110001", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            1167 => (0 => "01110000", 1 => "01110001", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            1168 => (0 => "11110010", 1 => "01110010", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            1169 => (0 => "00110010", 1 => "01110010", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            1170 => (0 => "01010010", 1 => "01110010", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            1171 => (0 => "01100010", 1 => "01110010", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            1172 => (0 => "01111010", 1 => "01110010", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            1173 => (0 => "01110110", 1 => "01110010", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            1174 => (0 => "01110000", 1 => "01110010", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            1175 => (0 => "01110011", 1 => "01110010", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            1176 => (0 => "11110011", 1 => "01110011", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            1177 => (0 => "00110011", 1 => "01110011", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            1178 => (0 => "01010011", 1 => "01110011", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            1179 => (0 => "01100011", 1 => "01110011", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            1180 => (0 => "01111011", 1 => "01110011", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            1181 => (0 => "01110111", 1 => "01110011", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            1182 => (0 => "01110001", 1 => "01110011", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            1183 => (0 => "01110010", 1 => "01110011", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            1184 => (0 => "11110100", 1 => "01110100", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            1185 => (0 => "00110100", 1 => "01110100", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            1186 => (0 => "01010100", 1 => "01110100", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            1187 => (0 => "01100100", 1 => "01110100", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            1188 => (0 => "01111100", 1 => "01110100", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            1189 => (0 => "01110000", 1 => "01110100", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            1190 => (0 => "01110110", 1 => "01110100", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            1191 => (0 => "01110101", 1 => "01110100", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            1192 => (0 => "11110101", 1 => "01110101", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            1193 => (0 => "00110101", 1 => "01110101", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            1194 => (0 => "01010101", 1 => "01110101", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            1195 => (0 => "01100101", 1 => "01110101", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            1196 => (0 => "01111101", 1 => "01110101", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            1197 => (0 => "01110001", 1 => "01110101", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            1198 => (0 => "01110111", 1 => "01110101", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            1199 => (0 => "01110100", 1 => "01110101", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            1200 => (0 => "11110110", 1 => "01110110", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            1201 => (0 => "00110110", 1 => "01110110", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            1202 => (0 => "01010110", 1 => "01110110", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            1203 => (0 => "01100110", 1 => "01110110", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            1204 => (0 => "01111110", 1 => "01110110", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            1205 => (0 => "01110010", 1 => "01110110", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            1206 => (0 => "01110100", 1 => "01110110", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            1207 => (0 => "01110111", 1 => "01110110", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            1208 => (0 => "11110111", 1 => "01110111", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            1209 => (0 => "00110111", 1 => "01110111", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            1210 => (0 => "01010111", 1 => "01110111", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            1211 => (0 => "01100111", 1 => "01110111", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            1212 => (0 => "01111111", 1 => "01110111", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            1213 => (0 => "01110011", 1 => "01110111", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            1214 => (0 => "01110101", 1 => "01110111", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            1215 => (0 => "01110110", 1 => "01110111", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            1216 => (0 => "11111000", 1 => "01111000", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            1217 => (0 => "00111000", 1 => "01111000", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            1218 => (0 => "01011000", 1 => "01111000", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            1219 => (0 => "01101000", 1 => "01111000", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            1220 => (0 => "01110000", 1 => "01111000", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            1221 => (0 => "01111100", 1 => "01111000", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            1222 => (0 => "01111010", 1 => "01111000", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            1223 => (0 => "01111001", 1 => "01111000", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            1224 => (0 => "11111001", 1 => "01111001", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            1225 => (0 => "00111001", 1 => "01111001", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            1226 => (0 => "01011001", 1 => "01111001", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            1227 => (0 => "01101001", 1 => "01111001", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            1228 => (0 => "01110001", 1 => "01111001", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            1229 => (0 => "01111101", 1 => "01111001", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            1230 => (0 => "01111011", 1 => "01111001", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            1231 => (0 => "01111000", 1 => "01111001", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            1232 => (0 => "11111010", 1 => "01111010", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            1233 => (0 => "00111010", 1 => "01111010", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            1234 => (0 => "01011010", 1 => "01111010", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            1235 => (0 => "01101010", 1 => "01111010", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            1236 => (0 => "01110010", 1 => "01111010", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            1237 => (0 => "01111110", 1 => "01111010", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            1238 => (0 => "01111000", 1 => "01111010", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            1239 => (0 => "01111011", 1 => "01111010", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            1240 => (0 => "11111011", 1 => "01111011", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            1241 => (0 => "00111011", 1 => "01111011", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            1242 => (0 => "01011011", 1 => "01111011", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            1243 => (0 => "01101011", 1 => "01111011", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            1244 => (0 => "01110011", 1 => "01111011", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            1245 => (0 => "01111111", 1 => "01111011", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            1246 => (0 => "01111001", 1 => "01111011", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            1247 => (0 => "01111010", 1 => "01111011", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            1248 => (0 => "11111100", 1 => "01111100", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            1249 => (0 => "00111100", 1 => "01111100", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            1250 => (0 => "01011100", 1 => "01111100", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            1251 => (0 => "01101100", 1 => "01111100", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            1252 => (0 => "01110100", 1 => "01111100", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            1253 => (0 => "01111000", 1 => "01111100", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            1254 => (0 => "01111110", 1 => "01111100", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            1255 => (0 => "01111101", 1 => "01111100", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            1256 => (0 => "11111101", 1 => "01111101", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            1257 => (0 => "00111101", 1 => "01111101", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            1258 => (0 => "01011101", 1 => "01111101", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            1259 => (0 => "01101101", 1 => "01111101", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            1260 => (0 => "01110101", 1 => "01111101", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            1261 => (0 => "01111001", 1 => "01111101", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            1262 => (0 => "01111111", 1 => "01111101", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            1263 => (0 => "01111100", 1 => "01111101", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            1264 => (0 => "11111110", 1 => "01111110", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            1265 => (0 => "00111110", 1 => "01111110", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            1266 => (0 => "01011110", 1 => "01111110", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            1267 => (0 => "01101110", 1 => "01111110", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            1268 => (0 => "01110110", 1 => "01111110", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            1269 => (0 => "01111010", 1 => "01111110", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            1270 => (0 => "01111100", 1 => "01111110", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            1271 => (0 => "01111111", 1 => "01111110", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            1272 => (0 => "11111111", 1 => "01111111", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            1273 => (0 => "00111111", 1 => "01111111", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            1274 => (0 => "01011111", 1 => "01111111", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            1275 => (0 => "01101111", 1 => "01111111", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            1276 => (0 => "01110111", 1 => "01111111", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            1277 => (0 => "01111011", 1 => "01111111", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            1278 => (0 => "01111101", 1 => "01111111", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            1279 => (0 => "01111110", 1 => "01111111", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            1280 => (0 => "00000000", 1 => "10000000", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            1281 => (0 => "11000000", 1 => "10000000", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            1282 => (0 => "10100000", 1 => "10000000", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            1283 => (0 => "10010000", 1 => "10000000", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            1284 => (0 => "10001000", 1 => "10000000", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            1285 => (0 => "10000100", 1 => "10000000", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            1286 => (0 => "10000010", 1 => "10000000", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            1287 => (0 => "10000001", 1 => "10000000", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            1288 => (0 => "00000001", 1 => "10000001", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            1289 => (0 => "11000001", 1 => "10000001", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            1290 => (0 => "10100001", 1 => "10000001", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            1291 => (0 => "10010001", 1 => "10000001", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            1292 => (0 => "10001001", 1 => "10000001", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            1293 => (0 => "10000101", 1 => "10000001", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            1294 => (0 => "10000011", 1 => "10000001", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            1295 => (0 => "10000000", 1 => "10000001", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            1296 => (0 => "00000010", 1 => "10000010", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            1297 => (0 => "11000010", 1 => "10000010", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            1298 => (0 => "10100010", 1 => "10000010", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            1299 => (0 => "10010010", 1 => "10000010", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            1300 => (0 => "10001010", 1 => "10000010", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            1301 => (0 => "10000110", 1 => "10000010", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            1302 => (0 => "10000000", 1 => "10000010", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            1303 => (0 => "10000011", 1 => "10000010", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            1304 => (0 => "00000011", 1 => "10000011", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            1305 => (0 => "11000011", 1 => "10000011", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            1306 => (0 => "10100011", 1 => "10000011", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            1307 => (0 => "10010011", 1 => "10000011", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            1308 => (0 => "10001011", 1 => "10000011", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            1309 => (0 => "10000111", 1 => "10000011", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            1310 => (0 => "10000001", 1 => "10000011", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            1311 => (0 => "10000010", 1 => "10000011", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            1312 => (0 => "00000100", 1 => "10000100", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            1313 => (0 => "11000100", 1 => "10000100", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            1314 => (0 => "10100100", 1 => "10000100", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            1315 => (0 => "10010100", 1 => "10000100", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            1316 => (0 => "10001100", 1 => "10000100", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            1317 => (0 => "10000000", 1 => "10000100", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            1318 => (0 => "10000110", 1 => "10000100", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            1319 => (0 => "10000101", 1 => "10000100", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            1320 => (0 => "00000101", 1 => "10000101", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            1321 => (0 => "11000101", 1 => "10000101", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            1322 => (0 => "10100101", 1 => "10000101", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            1323 => (0 => "10010101", 1 => "10000101", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            1324 => (0 => "10001101", 1 => "10000101", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            1325 => (0 => "10000001", 1 => "10000101", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            1326 => (0 => "10000111", 1 => "10000101", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            1327 => (0 => "10000100", 1 => "10000101", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            1328 => (0 => "00000110", 1 => "10000110", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            1329 => (0 => "11000110", 1 => "10000110", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            1330 => (0 => "10100110", 1 => "10000110", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            1331 => (0 => "10010110", 1 => "10000110", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            1332 => (0 => "10001110", 1 => "10000110", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            1333 => (0 => "10000010", 1 => "10000110", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            1334 => (0 => "10000100", 1 => "10000110", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            1335 => (0 => "10000111", 1 => "10000110", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            1336 => (0 => "00000111", 1 => "10000111", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            1337 => (0 => "11000111", 1 => "10000111", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            1338 => (0 => "10100111", 1 => "10000111", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            1339 => (0 => "10010111", 1 => "10000111", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            1340 => (0 => "10001111", 1 => "10000111", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            1341 => (0 => "10000011", 1 => "10000111", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            1342 => (0 => "10000101", 1 => "10000111", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            1343 => (0 => "10000110", 1 => "10000111", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            1344 => (0 => "00001000", 1 => "10001000", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            1345 => (0 => "11001000", 1 => "10001000", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            1346 => (0 => "10101000", 1 => "10001000", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            1347 => (0 => "10011000", 1 => "10001000", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            1348 => (0 => "10000000", 1 => "10001000", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            1349 => (0 => "10001100", 1 => "10001000", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            1350 => (0 => "10001010", 1 => "10001000", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            1351 => (0 => "10001001", 1 => "10001000", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            1352 => (0 => "00001001", 1 => "10001001", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            1353 => (0 => "11001001", 1 => "10001001", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            1354 => (0 => "10101001", 1 => "10001001", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            1355 => (0 => "10011001", 1 => "10001001", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            1356 => (0 => "10000001", 1 => "10001001", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            1357 => (0 => "10001101", 1 => "10001001", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            1358 => (0 => "10001011", 1 => "10001001", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            1359 => (0 => "10001000", 1 => "10001001", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            1360 => (0 => "00001010", 1 => "10001010", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            1361 => (0 => "11001010", 1 => "10001010", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            1362 => (0 => "10101010", 1 => "10001010", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            1363 => (0 => "10011010", 1 => "10001010", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            1364 => (0 => "10000010", 1 => "10001010", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            1365 => (0 => "10001110", 1 => "10001010", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            1366 => (0 => "10001000", 1 => "10001010", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            1367 => (0 => "10001011", 1 => "10001010", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            1368 => (0 => "00001011", 1 => "10001011", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            1369 => (0 => "11001011", 1 => "10001011", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            1370 => (0 => "10101011", 1 => "10001011", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            1371 => (0 => "10011011", 1 => "10001011", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            1372 => (0 => "10000011", 1 => "10001011", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            1373 => (0 => "10001111", 1 => "10001011", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            1374 => (0 => "10001001", 1 => "10001011", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            1375 => (0 => "10001010", 1 => "10001011", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            1376 => (0 => "00001100", 1 => "10001100", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            1377 => (0 => "11001100", 1 => "10001100", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            1378 => (0 => "10101100", 1 => "10001100", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            1379 => (0 => "10011100", 1 => "10001100", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            1380 => (0 => "10000100", 1 => "10001100", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            1381 => (0 => "10001000", 1 => "10001100", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            1382 => (0 => "10001110", 1 => "10001100", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            1383 => (0 => "10001101", 1 => "10001100", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            1384 => (0 => "00001101", 1 => "10001101", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            1385 => (0 => "11001101", 1 => "10001101", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            1386 => (0 => "10101101", 1 => "10001101", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            1387 => (0 => "10011101", 1 => "10001101", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            1388 => (0 => "10000101", 1 => "10001101", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            1389 => (0 => "10001001", 1 => "10001101", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            1390 => (0 => "10001111", 1 => "10001101", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            1391 => (0 => "10001100", 1 => "10001101", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            1392 => (0 => "00001110", 1 => "10001110", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            1393 => (0 => "11001110", 1 => "10001110", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            1394 => (0 => "10101110", 1 => "10001110", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            1395 => (0 => "10011110", 1 => "10001110", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            1396 => (0 => "10000110", 1 => "10001110", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            1397 => (0 => "10001010", 1 => "10001110", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            1398 => (0 => "10001100", 1 => "10001110", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            1399 => (0 => "10001111", 1 => "10001110", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            1400 => (0 => "00001111", 1 => "10001111", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            1401 => (0 => "11001111", 1 => "10001111", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            1402 => (0 => "10101111", 1 => "10001111", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            1403 => (0 => "10011111", 1 => "10001111", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            1404 => (0 => "10000111", 1 => "10001111", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            1405 => (0 => "10001011", 1 => "10001111", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            1406 => (0 => "10001101", 1 => "10001111", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            1407 => (0 => "10001110", 1 => "10001111", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            1408 => (0 => "00010000", 1 => "10010000", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            1409 => (0 => "11010000", 1 => "10010000", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            1410 => (0 => "10110000", 1 => "10010000", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            1411 => (0 => "10000000", 1 => "10010000", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            1412 => (0 => "10011000", 1 => "10010000", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            1413 => (0 => "10010100", 1 => "10010000", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            1414 => (0 => "10010010", 1 => "10010000", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            1415 => (0 => "10010001", 1 => "10010000", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            1416 => (0 => "00010001", 1 => "10010001", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            1417 => (0 => "11010001", 1 => "10010001", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            1418 => (0 => "10110001", 1 => "10010001", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            1419 => (0 => "10000001", 1 => "10010001", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            1420 => (0 => "10011001", 1 => "10010001", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            1421 => (0 => "10010101", 1 => "10010001", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            1422 => (0 => "10010011", 1 => "10010001", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            1423 => (0 => "10010000", 1 => "10010001", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            1424 => (0 => "00010010", 1 => "10010010", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            1425 => (0 => "11010010", 1 => "10010010", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            1426 => (0 => "10110010", 1 => "10010010", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            1427 => (0 => "10000010", 1 => "10010010", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            1428 => (0 => "10011010", 1 => "10010010", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            1429 => (0 => "10010110", 1 => "10010010", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            1430 => (0 => "10010000", 1 => "10010010", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            1431 => (0 => "10010011", 1 => "10010010", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            1432 => (0 => "00010011", 1 => "10010011", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            1433 => (0 => "11010011", 1 => "10010011", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            1434 => (0 => "10110011", 1 => "10010011", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            1435 => (0 => "10000011", 1 => "10010011", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            1436 => (0 => "10011011", 1 => "10010011", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            1437 => (0 => "10010111", 1 => "10010011", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            1438 => (0 => "10010001", 1 => "10010011", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            1439 => (0 => "10010010", 1 => "10010011", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            1440 => (0 => "00010100", 1 => "10010100", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            1441 => (0 => "11010100", 1 => "10010100", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            1442 => (0 => "10110100", 1 => "10010100", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            1443 => (0 => "10000100", 1 => "10010100", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            1444 => (0 => "10011100", 1 => "10010100", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            1445 => (0 => "10010000", 1 => "10010100", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            1446 => (0 => "10010110", 1 => "10010100", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            1447 => (0 => "10010101", 1 => "10010100", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            1448 => (0 => "00010101", 1 => "10010101", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            1449 => (0 => "11010101", 1 => "10010101", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            1450 => (0 => "10110101", 1 => "10010101", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            1451 => (0 => "10000101", 1 => "10010101", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            1452 => (0 => "10011101", 1 => "10010101", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            1453 => (0 => "10010001", 1 => "10010101", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            1454 => (0 => "10010111", 1 => "10010101", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            1455 => (0 => "10010100", 1 => "10010101", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            1456 => (0 => "00010110", 1 => "10010110", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            1457 => (0 => "11010110", 1 => "10010110", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            1458 => (0 => "10110110", 1 => "10010110", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            1459 => (0 => "10000110", 1 => "10010110", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            1460 => (0 => "10011110", 1 => "10010110", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            1461 => (0 => "10010010", 1 => "10010110", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            1462 => (0 => "10010100", 1 => "10010110", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            1463 => (0 => "10010111", 1 => "10010110", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            1464 => (0 => "00010111", 1 => "10010111", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            1465 => (0 => "11010111", 1 => "10010111", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            1466 => (0 => "10110111", 1 => "10010111", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            1467 => (0 => "10000111", 1 => "10010111", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            1468 => (0 => "10011111", 1 => "10010111", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            1469 => (0 => "10010011", 1 => "10010111", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            1470 => (0 => "10010101", 1 => "10010111", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            1471 => (0 => "10010110", 1 => "10010111", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            1472 => (0 => "00011000", 1 => "10011000", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            1473 => (0 => "11011000", 1 => "10011000", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            1474 => (0 => "10111000", 1 => "10011000", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            1475 => (0 => "10001000", 1 => "10011000", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            1476 => (0 => "10010000", 1 => "10011000", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            1477 => (0 => "10011100", 1 => "10011000", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            1478 => (0 => "10011010", 1 => "10011000", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            1479 => (0 => "10011001", 1 => "10011000", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            1480 => (0 => "00011001", 1 => "10011001", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            1481 => (0 => "11011001", 1 => "10011001", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            1482 => (0 => "10111001", 1 => "10011001", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            1483 => (0 => "10001001", 1 => "10011001", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            1484 => (0 => "10010001", 1 => "10011001", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            1485 => (0 => "10011101", 1 => "10011001", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            1486 => (0 => "10011011", 1 => "10011001", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            1487 => (0 => "10011000", 1 => "10011001", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            1488 => (0 => "00011010", 1 => "10011010", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            1489 => (0 => "11011010", 1 => "10011010", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            1490 => (0 => "10111010", 1 => "10011010", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            1491 => (0 => "10001010", 1 => "10011010", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            1492 => (0 => "10010010", 1 => "10011010", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            1493 => (0 => "10011110", 1 => "10011010", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            1494 => (0 => "10011000", 1 => "10011010", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            1495 => (0 => "10011011", 1 => "10011010", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            1496 => (0 => "00011011", 1 => "10011011", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            1497 => (0 => "11011011", 1 => "10011011", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            1498 => (0 => "10111011", 1 => "10011011", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            1499 => (0 => "10001011", 1 => "10011011", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            1500 => (0 => "10010011", 1 => "10011011", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            1501 => (0 => "10011111", 1 => "10011011", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            1502 => (0 => "10011001", 1 => "10011011", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            1503 => (0 => "10011010", 1 => "10011011", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            1504 => (0 => "00011100", 1 => "10011100", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            1505 => (0 => "11011100", 1 => "10011100", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            1506 => (0 => "10111100", 1 => "10011100", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            1507 => (0 => "10001100", 1 => "10011100", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            1508 => (0 => "10010100", 1 => "10011100", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            1509 => (0 => "10011000", 1 => "10011100", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            1510 => (0 => "10011110", 1 => "10011100", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            1511 => (0 => "10011101", 1 => "10011100", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            1512 => (0 => "00011101", 1 => "10011101", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            1513 => (0 => "11011101", 1 => "10011101", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            1514 => (0 => "10111101", 1 => "10011101", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            1515 => (0 => "10001101", 1 => "10011101", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            1516 => (0 => "10010101", 1 => "10011101", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            1517 => (0 => "10011001", 1 => "10011101", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            1518 => (0 => "10011111", 1 => "10011101", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            1519 => (0 => "10011100", 1 => "10011101", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            1520 => (0 => "00011110", 1 => "10011110", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            1521 => (0 => "11011110", 1 => "10011110", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            1522 => (0 => "10111110", 1 => "10011110", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            1523 => (0 => "10001110", 1 => "10011110", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            1524 => (0 => "10010110", 1 => "10011110", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            1525 => (0 => "10011010", 1 => "10011110", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            1526 => (0 => "10011100", 1 => "10011110", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            1527 => (0 => "10011111", 1 => "10011110", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            1528 => (0 => "00011111", 1 => "10011111", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            1529 => (0 => "11011111", 1 => "10011111", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            1530 => (0 => "10111111", 1 => "10011111", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            1531 => (0 => "10001111", 1 => "10011111", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            1532 => (0 => "10010111", 1 => "10011111", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            1533 => (0 => "10011011", 1 => "10011111", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            1534 => (0 => "10011101", 1 => "10011111", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            1535 => (0 => "10011110", 1 => "10011111", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            1536 => (0 => "00100000", 1 => "10100000", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            1537 => (0 => "11100000", 1 => "10100000", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            1538 => (0 => "10000000", 1 => "10100000", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            1539 => (0 => "10110000", 1 => "10100000", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            1540 => (0 => "10101000", 1 => "10100000", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            1541 => (0 => "10100100", 1 => "10100000", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            1542 => (0 => "10100010", 1 => "10100000", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            1543 => (0 => "10100001", 1 => "10100000", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            1544 => (0 => "00100001", 1 => "10100001", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            1545 => (0 => "11100001", 1 => "10100001", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            1546 => (0 => "10000001", 1 => "10100001", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            1547 => (0 => "10110001", 1 => "10100001", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            1548 => (0 => "10101001", 1 => "10100001", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            1549 => (0 => "10100101", 1 => "10100001", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            1550 => (0 => "10100011", 1 => "10100001", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            1551 => (0 => "10100000", 1 => "10100001", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            1552 => (0 => "00100010", 1 => "10100010", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            1553 => (0 => "11100010", 1 => "10100010", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            1554 => (0 => "10000010", 1 => "10100010", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            1555 => (0 => "10110010", 1 => "10100010", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            1556 => (0 => "10101010", 1 => "10100010", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            1557 => (0 => "10100110", 1 => "10100010", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            1558 => (0 => "10100000", 1 => "10100010", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            1559 => (0 => "10100011", 1 => "10100010", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            1560 => (0 => "00100011", 1 => "10100011", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            1561 => (0 => "11100011", 1 => "10100011", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            1562 => (0 => "10000011", 1 => "10100011", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            1563 => (0 => "10110011", 1 => "10100011", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            1564 => (0 => "10101011", 1 => "10100011", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            1565 => (0 => "10100111", 1 => "10100011", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            1566 => (0 => "10100001", 1 => "10100011", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            1567 => (0 => "10100010", 1 => "10100011", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            1568 => (0 => "00100100", 1 => "10100100", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            1569 => (0 => "11100100", 1 => "10100100", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            1570 => (0 => "10000100", 1 => "10100100", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            1571 => (0 => "10110100", 1 => "10100100", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            1572 => (0 => "10101100", 1 => "10100100", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            1573 => (0 => "10100000", 1 => "10100100", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            1574 => (0 => "10100110", 1 => "10100100", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            1575 => (0 => "10100101", 1 => "10100100", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            1576 => (0 => "00100101", 1 => "10100101", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            1577 => (0 => "11100101", 1 => "10100101", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            1578 => (0 => "10000101", 1 => "10100101", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            1579 => (0 => "10110101", 1 => "10100101", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            1580 => (0 => "10101101", 1 => "10100101", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            1581 => (0 => "10100001", 1 => "10100101", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            1582 => (0 => "10100111", 1 => "10100101", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            1583 => (0 => "10100100", 1 => "10100101", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            1584 => (0 => "00100110", 1 => "10100110", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            1585 => (0 => "11100110", 1 => "10100110", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            1586 => (0 => "10000110", 1 => "10100110", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            1587 => (0 => "10110110", 1 => "10100110", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            1588 => (0 => "10101110", 1 => "10100110", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            1589 => (0 => "10100010", 1 => "10100110", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            1590 => (0 => "10100100", 1 => "10100110", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            1591 => (0 => "10100111", 1 => "10100110", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            1592 => (0 => "00100111", 1 => "10100111", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            1593 => (0 => "11100111", 1 => "10100111", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            1594 => (0 => "10000111", 1 => "10100111", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            1595 => (0 => "10110111", 1 => "10100111", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            1596 => (0 => "10101111", 1 => "10100111", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            1597 => (0 => "10100011", 1 => "10100111", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            1598 => (0 => "10100101", 1 => "10100111", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            1599 => (0 => "10100110", 1 => "10100111", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            1600 => (0 => "00101000", 1 => "10101000", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            1601 => (0 => "11101000", 1 => "10101000", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            1602 => (0 => "10001000", 1 => "10101000", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            1603 => (0 => "10111000", 1 => "10101000", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            1604 => (0 => "10100000", 1 => "10101000", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            1605 => (0 => "10101100", 1 => "10101000", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            1606 => (0 => "10101010", 1 => "10101000", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            1607 => (0 => "10101001", 1 => "10101000", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            1608 => (0 => "00101001", 1 => "10101001", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            1609 => (0 => "11101001", 1 => "10101001", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            1610 => (0 => "10001001", 1 => "10101001", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            1611 => (0 => "10111001", 1 => "10101001", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            1612 => (0 => "10100001", 1 => "10101001", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            1613 => (0 => "10101101", 1 => "10101001", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            1614 => (0 => "10101011", 1 => "10101001", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            1615 => (0 => "10101000", 1 => "10101001", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            1616 => (0 => "00101010", 1 => "10101010", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            1617 => (0 => "11101010", 1 => "10101010", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            1618 => (0 => "10001010", 1 => "10101010", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            1619 => (0 => "10111010", 1 => "10101010", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            1620 => (0 => "10100010", 1 => "10101010", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            1621 => (0 => "10101110", 1 => "10101010", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            1622 => (0 => "10101000", 1 => "10101010", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            1623 => (0 => "10101011", 1 => "10101010", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            1624 => (0 => "00101011", 1 => "10101011", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            1625 => (0 => "11101011", 1 => "10101011", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            1626 => (0 => "10001011", 1 => "10101011", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            1627 => (0 => "10111011", 1 => "10101011", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            1628 => (0 => "10100011", 1 => "10101011", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            1629 => (0 => "10101111", 1 => "10101011", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            1630 => (0 => "10101001", 1 => "10101011", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            1631 => (0 => "10101010", 1 => "10101011", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            1632 => (0 => "00101100", 1 => "10101100", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            1633 => (0 => "11101100", 1 => "10101100", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            1634 => (0 => "10001100", 1 => "10101100", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            1635 => (0 => "10111100", 1 => "10101100", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            1636 => (0 => "10100100", 1 => "10101100", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            1637 => (0 => "10101000", 1 => "10101100", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            1638 => (0 => "10101110", 1 => "10101100", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            1639 => (0 => "10101101", 1 => "10101100", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            1640 => (0 => "00101101", 1 => "10101101", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            1641 => (0 => "11101101", 1 => "10101101", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            1642 => (0 => "10001101", 1 => "10101101", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            1643 => (0 => "10111101", 1 => "10101101", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            1644 => (0 => "10100101", 1 => "10101101", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            1645 => (0 => "10101001", 1 => "10101101", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            1646 => (0 => "10101111", 1 => "10101101", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            1647 => (0 => "10101100", 1 => "10101101", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            1648 => (0 => "00101110", 1 => "10101110", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            1649 => (0 => "11101110", 1 => "10101110", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            1650 => (0 => "10001110", 1 => "10101110", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            1651 => (0 => "10111110", 1 => "10101110", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            1652 => (0 => "10100110", 1 => "10101110", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            1653 => (0 => "10101010", 1 => "10101110", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            1654 => (0 => "10101100", 1 => "10101110", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            1655 => (0 => "10101111", 1 => "10101110", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            1656 => (0 => "00101111", 1 => "10101111", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            1657 => (0 => "11101111", 1 => "10101111", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            1658 => (0 => "10001111", 1 => "10101111", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            1659 => (0 => "10111111", 1 => "10101111", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            1660 => (0 => "10100111", 1 => "10101111", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            1661 => (0 => "10101011", 1 => "10101111", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            1662 => (0 => "10101101", 1 => "10101111", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            1663 => (0 => "10101110", 1 => "10101111", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            1664 => (0 => "00110000", 1 => "10110000", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            1665 => (0 => "11110000", 1 => "10110000", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            1666 => (0 => "10010000", 1 => "10110000", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            1667 => (0 => "10100000", 1 => "10110000", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            1668 => (0 => "10111000", 1 => "10110000", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            1669 => (0 => "10110100", 1 => "10110000", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            1670 => (0 => "10110010", 1 => "10110000", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            1671 => (0 => "10110001", 1 => "10110000", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            1672 => (0 => "00110001", 1 => "10110001", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            1673 => (0 => "11110001", 1 => "10110001", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            1674 => (0 => "10010001", 1 => "10110001", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            1675 => (0 => "10100001", 1 => "10110001", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            1676 => (0 => "10111001", 1 => "10110001", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            1677 => (0 => "10110101", 1 => "10110001", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            1678 => (0 => "10110011", 1 => "10110001", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            1679 => (0 => "10110000", 1 => "10110001", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            1680 => (0 => "00110010", 1 => "10110010", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            1681 => (0 => "11110010", 1 => "10110010", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            1682 => (0 => "10010010", 1 => "10110010", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            1683 => (0 => "10100010", 1 => "10110010", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            1684 => (0 => "10111010", 1 => "10110010", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            1685 => (0 => "10110110", 1 => "10110010", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            1686 => (0 => "10110000", 1 => "10110010", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            1687 => (0 => "10110011", 1 => "10110010", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            1688 => (0 => "00110011", 1 => "10110011", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            1689 => (0 => "11110011", 1 => "10110011", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            1690 => (0 => "10010011", 1 => "10110011", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            1691 => (0 => "10100011", 1 => "10110011", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            1692 => (0 => "10111011", 1 => "10110011", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            1693 => (0 => "10110111", 1 => "10110011", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            1694 => (0 => "10110001", 1 => "10110011", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            1695 => (0 => "10110010", 1 => "10110011", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            1696 => (0 => "00110100", 1 => "10110100", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            1697 => (0 => "11110100", 1 => "10110100", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            1698 => (0 => "10010100", 1 => "10110100", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            1699 => (0 => "10100100", 1 => "10110100", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            1700 => (0 => "10111100", 1 => "10110100", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            1701 => (0 => "10110000", 1 => "10110100", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            1702 => (0 => "10110110", 1 => "10110100", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            1703 => (0 => "10110101", 1 => "10110100", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            1704 => (0 => "00110101", 1 => "10110101", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            1705 => (0 => "11110101", 1 => "10110101", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            1706 => (0 => "10010101", 1 => "10110101", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            1707 => (0 => "10100101", 1 => "10110101", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            1708 => (0 => "10111101", 1 => "10110101", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            1709 => (0 => "10110001", 1 => "10110101", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            1710 => (0 => "10110111", 1 => "10110101", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            1711 => (0 => "10110100", 1 => "10110101", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            1712 => (0 => "00110110", 1 => "10110110", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            1713 => (0 => "11110110", 1 => "10110110", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            1714 => (0 => "10010110", 1 => "10110110", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            1715 => (0 => "10100110", 1 => "10110110", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            1716 => (0 => "10111110", 1 => "10110110", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            1717 => (0 => "10110010", 1 => "10110110", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            1718 => (0 => "10110100", 1 => "10110110", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            1719 => (0 => "10110111", 1 => "10110110", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            1720 => (0 => "00110111", 1 => "10110111", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            1721 => (0 => "11110111", 1 => "10110111", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            1722 => (0 => "10010111", 1 => "10110111", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            1723 => (0 => "10100111", 1 => "10110111", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            1724 => (0 => "10111111", 1 => "10110111", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            1725 => (0 => "10110011", 1 => "10110111", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            1726 => (0 => "10110101", 1 => "10110111", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            1727 => (0 => "10110110", 1 => "10110111", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            1728 => (0 => "00111000", 1 => "10111000", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            1729 => (0 => "11111000", 1 => "10111000", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            1730 => (0 => "10011000", 1 => "10111000", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            1731 => (0 => "10101000", 1 => "10111000", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            1732 => (0 => "10110000", 1 => "10111000", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            1733 => (0 => "10111100", 1 => "10111000", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            1734 => (0 => "10111010", 1 => "10111000", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            1735 => (0 => "10111001", 1 => "10111000", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            1736 => (0 => "00111001", 1 => "10111001", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            1737 => (0 => "11111001", 1 => "10111001", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            1738 => (0 => "10011001", 1 => "10111001", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            1739 => (0 => "10101001", 1 => "10111001", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            1740 => (0 => "10110001", 1 => "10111001", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            1741 => (0 => "10111101", 1 => "10111001", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            1742 => (0 => "10111011", 1 => "10111001", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            1743 => (0 => "10111000", 1 => "10111001", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            1744 => (0 => "00111010", 1 => "10111010", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            1745 => (0 => "11111010", 1 => "10111010", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            1746 => (0 => "10011010", 1 => "10111010", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            1747 => (0 => "10101010", 1 => "10111010", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            1748 => (0 => "10110010", 1 => "10111010", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            1749 => (0 => "10111110", 1 => "10111010", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            1750 => (0 => "10111000", 1 => "10111010", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            1751 => (0 => "10111011", 1 => "10111010", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            1752 => (0 => "00111011", 1 => "10111011", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            1753 => (0 => "11111011", 1 => "10111011", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            1754 => (0 => "10011011", 1 => "10111011", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            1755 => (0 => "10101011", 1 => "10111011", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            1756 => (0 => "10110011", 1 => "10111011", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            1757 => (0 => "10111111", 1 => "10111011", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            1758 => (0 => "10111001", 1 => "10111011", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            1759 => (0 => "10111010", 1 => "10111011", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            1760 => (0 => "00111100", 1 => "10111100", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            1761 => (0 => "11111100", 1 => "10111100", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            1762 => (0 => "10011100", 1 => "10111100", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            1763 => (0 => "10101100", 1 => "10111100", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            1764 => (0 => "10110100", 1 => "10111100", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            1765 => (0 => "10111000", 1 => "10111100", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            1766 => (0 => "10111110", 1 => "10111100", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            1767 => (0 => "10111101", 1 => "10111100", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            1768 => (0 => "00111101", 1 => "10111101", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            1769 => (0 => "11111101", 1 => "10111101", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            1770 => (0 => "10011101", 1 => "10111101", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            1771 => (0 => "10101101", 1 => "10111101", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            1772 => (0 => "10110101", 1 => "10111101", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            1773 => (0 => "10111001", 1 => "10111101", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            1774 => (0 => "10111111", 1 => "10111101", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            1775 => (0 => "10111100", 1 => "10111101", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            1776 => (0 => "00111110", 1 => "10111110", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            1777 => (0 => "11111110", 1 => "10111110", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            1778 => (0 => "10011110", 1 => "10111110", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            1779 => (0 => "10101110", 1 => "10111110", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            1780 => (0 => "10110110", 1 => "10111110", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            1781 => (0 => "10111010", 1 => "10111110", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            1782 => (0 => "10111100", 1 => "10111110", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            1783 => (0 => "10111111", 1 => "10111110", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            1784 => (0 => "00111111", 1 => "10111111", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            1785 => (0 => "11111111", 1 => "10111111", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            1786 => (0 => "10011111", 1 => "10111111", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            1787 => (0 => "10101111", 1 => "10111111", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            1788 => (0 => "10110111", 1 => "10111111", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            1789 => (0 => "10111011", 1 => "10111111", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            1790 => (0 => "10111101", 1 => "10111111", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            1791 => (0 => "10111110", 1 => "10111111", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            1792 => (0 => "01000000", 1 => "11000000", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            1793 => (0 => "10000000", 1 => "11000000", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            1794 => (0 => "11100000", 1 => "11000000", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            1795 => (0 => "11010000", 1 => "11000000", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            1796 => (0 => "11001000", 1 => "11000000", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            1797 => (0 => "11000100", 1 => "11000000", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            1798 => (0 => "11000010", 1 => "11000000", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            1799 => (0 => "11000001", 1 => "11000000", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            1800 => (0 => "01000001", 1 => "11000001", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            1801 => (0 => "10000001", 1 => "11000001", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            1802 => (0 => "11100001", 1 => "11000001", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            1803 => (0 => "11010001", 1 => "11000001", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            1804 => (0 => "11001001", 1 => "11000001", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            1805 => (0 => "11000101", 1 => "11000001", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            1806 => (0 => "11000011", 1 => "11000001", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            1807 => (0 => "11000000", 1 => "11000001", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            1808 => (0 => "01000010", 1 => "11000010", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            1809 => (0 => "10000010", 1 => "11000010", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            1810 => (0 => "11100010", 1 => "11000010", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            1811 => (0 => "11010010", 1 => "11000010", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            1812 => (0 => "11001010", 1 => "11000010", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            1813 => (0 => "11000110", 1 => "11000010", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            1814 => (0 => "11000000", 1 => "11000010", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            1815 => (0 => "11000011", 1 => "11000010", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            1816 => (0 => "01000011", 1 => "11000011", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            1817 => (0 => "10000011", 1 => "11000011", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            1818 => (0 => "11100011", 1 => "11000011", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            1819 => (0 => "11010011", 1 => "11000011", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            1820 => (0 => "11001011", 1 => "11000011", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            1821 => (0 => "11000111", 1 => "11000011", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            1822 => (0 => "11000001", 1 => "11000011", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            1823 => (0 => "11000010", 1 => "11000011", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            1824 => (0 => "01000100", 1 => "11000100", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            1825 => (0 => "10000100", 1 => "11000100", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            1826 => (0 => "11100100", 1 => "11000100", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            1827 => (0 => "11010100", 1 => "11000100", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            1828 => (0 => "11001100", 1 => "11000100", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            1829 => (0 => "11000000", 1 => "11000100", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            1830 => (0 => "11000110", 1 => "11000100", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            1831 => (0 => "11000101", 1 => "11000100", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            1832 => (0 => "01000101", 1 => "11000101", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            1833 => (0 => "10000101", 1 => "11000101", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            1834 => (0 => "11100101", 1 => "11000101", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            1835 => (0 => "11010101", 1 => "11000101", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            1836 => (0 => "11001101", 1 => "11000101", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            1837 => (0 => "11000001", 1 => "11000101", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            1838 => (0 => "11000111", 1 => "11000101", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            1839 => (0 => "11000100", 1 => "11000101", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            1840 => (0 => "01000110", 1 => "11000110", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            1841 => (0 => "10000110", 1 => "11000110", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            1842 => (0 => "11100110", 1 => "11000110", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            1843 => (0 => "11010110", 1 => "11000110", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            1844 => (0 => "11001110", 1 => "11000110", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            1845 => (0 => "11000010", 1 => "11000110", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            1846 => (0 => "11000100", 1 => "11000110", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            1847 => (0 => "11000111", 1 => "11000110", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            1848 => (0 => "01000111", 1 => "11000111", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            1849 => (0 => "10000111", 1 => "11000111", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            1850 => (0 => "11100111", 1 => "11000111", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            1851 => (0 => "11010111", 1 => "11000111", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            1852 => (0 => "11001111", 1 => "11000111", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            1853 => (0 => "11000011", 1 => "11000111", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            1854 => (0 => "11000101", 1 => "11000111", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            1855 => (0 => "11000110", 1 => "11000111", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            1856 => (0 => "01001000", 1 => "11001000", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            1857 => (0 => "10001000", 1 => "11001000", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            1858 => (0 => "11101000", 1 => "11001000", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            1859 => (0 => "11011000", 1 => "11001000", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            1860 => (0 => "11000000", 1 => "11001000", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            1861 => (0 => "11001100", 1 => "11001000", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            1862 => (0 => "11001010", 1 => "11001000", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            1863 => (0 => "11001001", 1 => "11001000", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            1864 => (0 => "01001001", 1 => "11001001", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            1865 => (0 => "10001001", 1 => "11001001", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            1866 => (0 => "11101001", 1 => "11001001", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            1867 => (0 => "11011001", 1 => "11001001", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            1868 => (0 => "11000001", 1 => "11001001", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            1869 => (0 => "11001101", 1 => "11001001", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            1870 => (0 => "11001011", 1 => "11001001", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            1871 => (0 => "11001000", 1 => "11001001", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            1872 => (0 => "01001010", 1 => "11001010", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            1873 => (0 => "10001010", 1 => "11001010", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            1874 => (0 => "11101010", 1 => "11001010", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            1875 => (0 => "11011010", 1 => "11001010", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            1876 => (0 => "11000010", 1 => "11001010", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            1877 => (0 => "11001110", 1 => "11001010", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            1878 => (0 => "11001000", 1 => "11001010", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            1879 => (0 => "11001011", 1 => "11001010", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            1880 => (0 => "01001011", 1 => "11001011", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            1881 => (0 => "10001011", 1 => "11001011", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            1882 => (0 => "11101011", 1 => "11001011", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            1883 => (0 => "11011011", 1 => "11001011", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            1884 => (0 => "11000011", 1 => "11001011", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            1885 => (0 => "11001111", 1 => "11001011", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            1886 => (0 => "11001001", 1 => "11001011", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            1887 => (0 => "11001010", 1 => "11001011", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            1888 => (0 => "01001100", 1 => "11001100", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            1889 => (0 => "10001100", 1 => "11001100", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            1890 => (0 => "11101100", 1 => "11001100", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            1891 => (0 => "11011100", 1 => "11001100", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            1892 => (0 => "11000100", 1 => "11001100", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            1893 => (0 => "11001000", 1 => "11001100", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            1894 => (0 => "11001110", 1 => "11001100", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            1895 => (0 => "11001101", 1 => "11001100", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            1896 => (0 => "01001101", 1 => "11001101", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            1897 => (0 => "10001101", 1 => "11001101", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            1898 => (0 => "11101101", 1 => "11001101", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            1899 => (0 => "11011101", 1 => "11001101", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            1900 => (0 => "11000101", 1 => "11001101", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            1901 => (0 => "11001001", 1 => "11001101", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            1902 => (0 => "11001111", 1 => "11001101", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            1903 => (0 => "11001100", 1 => "11001101", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            1904 => (0 => "01001110", 1 => "11001110", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            1905 => (0 => "10001110", 1 => "11001110", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            1906 => (0 => "11101110", 1 => "11001110", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            1907 => (0 => "11011110", 1 => "11001110", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            1908 => (0 => "11000110", 1 => "11001110", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            1909 => (0 => "11001010", 1 => "11001110", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            1910 => (0 => "11001100", 1 => "11001110", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            1911 => (0 => "11001111", 1 => "11001110", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            1912 => (0 => "01001111", 1 => "11001111", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            1913 => (0 => "10001111", 1 => "11001111", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            1914 => (0 => "11101111", 1 => "11001111", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            1915 => (0 => "11011111", 1 => "11001111", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            1916 => (0 => "11000111", 1 => "11001111", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            1917 => (0 => "11001011", 1 => "11001111", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            1918 => (0 => "11001101", 1 => "11001111", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            1919 => (0 => "11001110", 1 => "11001111", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            1920 => (0 => "01010000", 1 => "11010000", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            1921 => (0 => "10010000", 1 => "11010000", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            1922 => (0 => "11110000", 1 => "11010000", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            1923 => (0 => "11000000", 1 => "11010000", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            1924 => (0 => "11011000", 1 => "11010000", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            1925 => (0 => "11010100", 1 => "11010000", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            1926 => (0 => "11010010", 1 => "11010000", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            1927 => (0 => "11010001", 1 => "11010000", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            1928 => (0 => "01010001", 1 => "11010001", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            1929 => (0 => "10010001", 1 => "11010001", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            1930 => (0 => "11110001", 1 => "11010001", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            1931 => (0 => "11000001", 1 => "11010001", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            1932 => (0 => "11011001", 1 => "11010001", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            1933 => (0 => "11010101", 1 => "11010001", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            1934 => (0 => "11010011", 1 => "11010001", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            1935 => (0 => "11010000", 1 => "11010001", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            1936 => (0 => "01010010", 1 => "11010010", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            1937 => (0 => "10010010", 1 => "11010010", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            1938 => (0 => "11110010", 1 => "11010010", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            1939 => (0 => "11000010", 1 => "11010010", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            1940 => (0 => "11011010", 1 => "11010010", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            1941 => (0 => "11010110", 1 => "11010010", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            1942 => (0 => "11010000", 1 => "11010010", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            1943 => (0 => "11010011", 1 => "11010010", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            1944 => (0 => "01010011", 1 => "11010011", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            1945 => (0 => "10010011", 1 => "11010011", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            1946 => (0 => "11110011", 1 => "11010011", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            1947 => (0 => "11000011", 1 => "11010011", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            1948 => (0 => "11011011", 1 => "11010011", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            1949 => (0 => "11010111", 1 => "11010011", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            1950 => (0 => "11010001", 1 => "11010011", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            1951 => (0 => "11010010", 1 => "11010011", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            1952 => (0 => "01010100", 1 => "11010100", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            1953 => (0 => "10010100", 1 => "11010100", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            1954 => (0 => "11110100", 1 => "11010100", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            1955 => (0 => "11000100", 1 => "11010100", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            1956 => (0 => "11011100", 1 => "11010100", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            1957 => (0 => "11010000", 1 => "11010100", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            1958 => (0 => "11010110", 1 => "11010100", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            1959 => (0 => "11010101", 1 => "11010100", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            1960 => (0 => "01010101", 1 => "11010101", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            1961 => (0 => "10010101", 1 => "11010101", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            1962 => (0 => "11110101", 1 => "11010101", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            1963 => (0 => "11000101", 1 => "11010101", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            1964 => (0 => "11011101", 1 => "11010101", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            1965 => (0 => "11010001", 1 => "11010101", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            1966 => (0 => "11010111", 1 => "11010101", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            1967 => (0 => "11010100", 1 => "11010101", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            1968 => (0 => "01010110", 1 => "11010110", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            1969 => (0 => "10010110", 1 => "11010110", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            1970 => (0 => "11110110", 1 => "11010110", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            1971 => (0 => "11000110", 1 => "11010110", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            1972 => (0 => "11011110", 1 => "11010110", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            1973 => (0 => "11010010", 1 => "11010110", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            1974 => (0 => "11010100", 1 => "11010110", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            1975 => (0 => "11010111", 1 => "11010110", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            1976 => (0 => "01010111", 1 => "11010111", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            1977 => (0 => "10010111", 1 => "11010111", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            1978 => (0 => "11110111", 1 => "11010111", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            1979 => (0 => "11000111", 1 => "11010111", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            1980 => (0 => "11011111", 1 => "11010111", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            1981 => (0 => "11010011", 1 => "11010111", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            1982 => (0 => "11010101", 1 => "11010111", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            1983 => (0 => "11010110", 1 => "11010111", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            1984 => (0 => "01011000", 1 => "11011000", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            1985 => (0 => "10011000", 1 => "11011000", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            1986 => (0 => "11111000", 1 => "11011000", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            1987 => (0 => "11001000", 1 => "11011000", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            1988 => (0 => "11010000", 1 => "11011000", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            1989 => (0 => "11011100", 1 => "11011000", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            1990 => (0 => "11011010", 1 => "11011000", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            1991 => (0 => "11011001", 1 => "11011000", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            1992 => (0 => "01011001", 1 => "11011001", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            1993 => (0 => "10011001", 1 => "11011001", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            1994 => (0 => "11111001", 1 => "11011001", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            1995 => (0 => "11001001", 1 => "11011001", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            1996 => (0 => "11010001", 1 => "11011001", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            1997 => (0 => "11011101", 1 => "11011001", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            1998 => (0 => "11011011", 1 => "11011001", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            1999 => (0 => "11011000", 1 => "11011001", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            2000 => (0 => "01011010", 1 => "11011010", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            2001 => (0 => "10011010", 1 => "11011010", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            2002 => (0 => "11111010", 1 => "11011010", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            2003 => (0 => "11001010", 1 => "11011010", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            2004 => (0 => "11010010", 1 => "11011010", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            2005 => (0 => "11011110", 1 => "11011010", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            2006 => (0 => "11011000", 1 => "11011010", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            2007 => (0 => "11011011", 1 => "11011010", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            2008 => (0 => "01011011", 1 => "11011011", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            2009 => (0 => "10011011", 1 => "11011011", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            2010 => (0 => "11111011", 1 => "11011011", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            2011 => (0 => "11001011", 1 => "11011011", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            2012 => (0 => "11010011", 1 => "11011011", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            2013 => (0 => "11011111", 1 => "11011011", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            2014 => (0 => "11011001", 1 => "11011011", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            2015 => (0 => "11011010", 1 => "11011011", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            2016 => (0 => "01011100", 1 => "11011100", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            2017 => (0 => "10011100", 1 => "11011100", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            2018 => (0 => "11111100", 1 => "11011100", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            2019 => (0 => "11001100", 1 => "11011100", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            2020 => (0 => "11010100", 1 => "11011100", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            2021 => (0 => "11011000", 1 => "11011100", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            2022 => (0 => "11011110", 1 => "11011100", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            2023 => (0 => "11011101", 1 => "11011100", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            2024 => (0 => "01011101", 1 => "11011101", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            2025 => (0 => "10011101", 1 => "11011101", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            2026 => (0 => "11111101", 1 => "11011101", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            2027 => (0 => "11001101", 1 => "11011101", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            2028 => (0 => "11010101", 1 => "11011101", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            2029 => (0 => "11011001", 1 => "11011101", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            2030 => (0 => "11011111", 1 => "11011101", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            2031 => (0 => "11011100", 1 => "11011101", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            2032 => (0 => "01011110", 1 => "11011110", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            2033 => (0 => "10011110", 1 => "11011110", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            2034 => (0 => "11111110", 1 => "11011110", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            2035 => (0 => "11001110", 1 => "11011110", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            2036 => (0 => "11010110", 1 => "11011110", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            2037 => (0 => "11011010", 1 => "11011110", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            2038 => (0 => "11011100", 1 => "11011110", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            2039 => (0 => "11011111", 1 => "11011110", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            2040 => (0 => "01011111", 1 => "11011111", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            2041 => (0 => "10011111", 1 => "11011111", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            2042 => (0 => "11111111", 1 => "11011111", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            2043 => (0 => "11001111", 1 => "11011111", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            2044 => (0 => "11010111", 1 => "11011111", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            2045 => (0 => "11011011", 1 => "11011111", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            2046 => (0 => "11011101", 1 => "11011111", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            2047 => (0 => "11011110", 1 => "11011111", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            2048 => (0 => "01100000", 1 => "11100000", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            2049 => (0 => "10100000", 1 => "11100000", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            2050 => (0 => "11000000", 1 => "11100000", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            2051 => (0 => "11110000", 1 => "11100000", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            2052 => (0 => "11101000", 1 => "11100000", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            2053 => (0 => "11100100", 1 => "11100000", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            2054 => (0 => "11100010", 1 => "11100000", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            2055 => (0 => "11100001", 1 => "11100000", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            2056 => (0 => "01100001", 1 => "11100001", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            2057 => (0 => "10100001", 1 => "11100001", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            2058 => (0 => "11000001", 1 => "11100001", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            2059 => (0 => "11110001", 1 => "11100001", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            2060 => (0 => "11101001", 1 => "11100001", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            2061 => (0 => "11100101", 1 => "11100001", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            2062 => (0 => "11100011", 1 => "11100001", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            2063 => (0 => "11100000", 1 => "11100001", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            2064 => (0 => "01100010", 1 => "11100010", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            2065 => (0 => "10100010", 1 => "11100010", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            2066 => (0 => "11000010", 1 => "11100010", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            2067 => (0 => "11110010", 1 => "11100010", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            2068 => (0 => "11101010", 1 => "11100010", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            2069 => (0 => "11100110", 1 => "11100010", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            2070 => (0 => "11100000", 1 => "11100010", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            2071 => (0 => "11100011", 1 => "11100010", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            2072 => (0 => "01100011", 1 => "11100011", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            2073 => (0 => "10100011", 1 => "11100011", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            2074 => (0 => "11000011", 1 => "11100011", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            2075 => (0 => "11110011", 1 => "11100011", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            2076 => (0 => "11101011", 1 => "11100011", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            2077 => (0 => "11100111", 1 => "11100011", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            2078 => (0 => "11100001", 1 => "11100011", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            2079 => (0 => "11100010", 1 => "11100011", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            2080 => (0 => "01100100", 1 => "11100100", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            2081 => (0 => "10100100", 1 => "11100100", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            2082 => (0 => "11000100", 1 => "11100100", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            2083 => (0 => "11110100", 1 => "11100100", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            2084 => (0 => "11101100", 1 => "11100100", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            2085 => (0 => "11100000", 1 => "11100100", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            2086 => (0 => "11100110", 1 => "11100100", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            2087 => (0 => "11100101", 1 => "11100100", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            2088 => (0 => "01100101", 1 => "11100101", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            2089 => (0 => "10100101", 1 => "11100101", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            2090 => (0 => "11000101", 1 => "11100101", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            2091 => (0 => "11110101", 1 => "11100101", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            2092 => (0 => "11101101", 1 => "11100101", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            2093 => (0 => "11100001", 1 => "11100101", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            2094 => (0 => "11100111", 1 => "11100101", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            2095 => (0 => "11100100", 1 => "11100101", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            2096 => (0 => "01100110", 1 => "11100110", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            2097 => (0 => "10100110", 1 => "11100110", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            2098 => (0 => "11000110", 1 => "11100110", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            2099 => (0 => "11110110", 1 => "11100110", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            2100 => (0 => "11101110", 1 => "11100110", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            2101 => (0 => "11100010", 1 => "11100110", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            2102 => (0 => "11100100", 1 => "11100110", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            2103 => (0 => "11100111", 1 => "11100110", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            2104 => (0 => "01100111", 1 => "11100111", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            2105 => (0 => "10100111", 1 => "11100111", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            2106 => (0 => "11000111", 1 => "11100111", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            2107 => (0 => "11110111", 1 => "11100111", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            2108 => (0 => "11101111", 1 => "11100111", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            2109 => (0 => "11100011", 1 => "11100111", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            2110 => (0 => "11100101", 1 => "11100111", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            2111 => (0 => "11100110", 1 => "11100111", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            2112 => (0 => "01101000", 1 => "11101000", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            2113 => (0 => "10101000", 1 => "11101000", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            2114 => (0 => "11001000", 1 => "11101000", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            2115 => (0 => "11111000", 1 => "11101000", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            2116 => (0 => "11100000", 1 => "11101000", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            2117 => (0 => "11101100", 1 => "11101000", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            2118 => (0 => "11101010", 1 => "11101000", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            2119 => (0 => "11101001", 1 => "11101000", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            2120 => (0 => "01101001", 1 => "11101001", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            2121 => (0 => "10101001", 1 => "11101001", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            2122 => (0 => "11001001", 1 => "11101001", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            2123 => (0 => "11111001", 1 => "11101001", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            2124 => (0 => "11100001", 1 => "11101001", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            2125 => (0 => "11101101", 1 => "11101001", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            2126 => (0 => "11101011", 1 => "11101001", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            2127 => (0 => "11101000", 1 => "11101001", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            2128 => (0 => "01101010", 1 => "11101010", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            2129 => (0 => "10101010", 1 => "11101010", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            2130 => (0 => "11001010", 1 => "11101010", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            2131 => (0 => "11111010", 1 => "11101010", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            2132 => (0 => "11100010", 1 => "11101010", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            2133 => (0 => "11101110", 1 => "11101010", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            2134 => (0 => "11101000", 1 => "11101010", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            2135 => (0 => "11101011", 1 => "11101010", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            2136 => (0 => "01101011", 1 => "11101011", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            2137 => (0 => "10101011", 1 => "11101011", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            2138 => (0 => "11001011", 1 => "11101011", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            2139 => (0 => "11111011", 1 => "11101011", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            2140 => (0 => "11100011", 1 => "11101011", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            2141 => (0 => "11101111", 1 => "11101011", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            2142 => (0 => "11101001", 1 => "11101011", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            2143 => (0 => "11101010", 1 => "11101011", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            2144 => (0 => "01101100", 1 => "11101100", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            2145 => (0 => "10101100", 1 => "11101100", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            2146 => (0 => "11001100", 1 => "11101100", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            2147 => (0 => "11111100", 1 => "11101100", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            2148 => (0 => "11100100", 1 => "11101100", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            2149 => (0 => "11101000", 1 => "11101100", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            2150 => (0 => "11101110", 1 => "11101100", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            2151 => (0 => "11101101", 1 => "11101100", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            2152 => (0 => "01101101", 1 => "11101101", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            2153 => (0 => "10101101", 1 => "11101101", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            2154 => (0 => "11001101", 1 => "11101101", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            2155 => (0 => "11111101", 1 => "11101101", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            2156 => (0 => "11100101", 1 => "11101101", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            2157 => (0 => "11101001", 1 => "11101101", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            2158 => (0 => "11101111", 1 => "11101101", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            2159 => (0 => "11101100", 1 => "11101101", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            2160 => (0 => "01101110", 1 => "11101110", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            2161 => (0 => "10101110", 1 => "11101110", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            2162 => (0 => "11001110", 1 => "11101110", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            2163 => (0 => "11111110", 1 => "11101110", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            2164 => (0 => "11100110", 1 => "11101110", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            2165 => (0 => "11101010", 1 => "11101110", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            2166 => (0 => "11101100", 1 => "11101110", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            2167 => (0 => "11101111", 1 => "11101110", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            2168 => (0 => "01101111", 1 => "11101111", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            2169 => (0 => "10101111", 1 => "11101111", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            2170 => (0 => "11001111", 1 => "11101111", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            2171 => (0 => "11111111", 1 => "11101111", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            2172 => (0 => "11100111", 1 => "11101111", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            2173 => (0 => "11101011", 1 => "11101111", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            2174 => (0 => "11101101", 1 => "11101111", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            2175 => (0 => "11101110", 1 => "11101111", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            2176 => (0 => "01110000", 1 => "11110000", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            2177 => (0 => "10110000", 1 => "11110000", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            2178 => (0 => "11010000", 1 => "11110000", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            2179 => (0 => "11100000", 1 => "11110000", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            2180 => (0 => "11111000", 1 => "11110000", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            2181 => (0 => "11110100", 1 => "11110000", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            2182 => (0 => "11110010", 1 => "11110000", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            2183 => (0 => "11110001", 1 => "11110000", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            2184 => (0 => "01110001", 1 => "11110001", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            2185 => (0 => "10110001", 1 => "11110001", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            2186 => (0 => "11010001", 1 => "11110001", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            2187 => (0 => "11100001", 1 => "11110001", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            2188 => (0 => "11111001", 1 => "11110001", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            2189 => (0 => "11110101", 1 => "11110001", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            2190 => (0 => "11110011", 1 => "11110001", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            2191 => (0 => "11110000", 1 => "11110001", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            2192 => (0 => "01110010", 1 => "11110010", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            2193 => (0 => "10110010", 1 => "11110010", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            2194 => (0 => "11010010", 1 => "11110010", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            2195 => (0 => "11100010", 1 => "11110010", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            2196 => (0 => "11111010", 1 => "11110010", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            2197 => (0 => "11110110", 1 => "11110010", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            2198 => (0 => "11110000", 1 => "11110010", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            2199 => (0 => "11110011", 1 => "11110010", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            2200 => (0 => "01110011", 1 => "11110011", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            2201 => (0 => "10110011", 1 => "11110011", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            2202 => (0 => "11010011", 1 => "11110011", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            2203 => (0 => "11100011", 1 => "11110011", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            2204 => (0 => "11111011", 1 => "11110011", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            2205 => (0 => "11110111", 1 => "11110011", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            2206 => (0 => "11110001", 1 => "11110011", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            2207 => (0 => "11110010", 1 => "11110011", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            2208 => (0 => "01110100", 1 => "11110100", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            2209 => (0 => "10110100", 1 => "11110100", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            2210 => (0 => "11010100", 1 => "11110100", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            2211 => (0 => "11100100", 1 => "11110100", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            2212 => (0 => "11111100", 1 => "11110100", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            2213 => (0 => "11110000", 1 => "11110100", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            2214 => (0 => "11110110", 1 => "11110100", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            2215 => (0 => "11110101", 1 => "11110100", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            2216 => (0 => "01110101", 1 => "11110101", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            2217 => (0 => "10110101", 1 => "11110101", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            2218 => (0 => "11010101", 1 => "11110101", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            2219 => (0 => "11100101", 1 => "11110101", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            2220 => (0 => "11111101", 1 => "11110101", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            2221 => (0 => "11110001", 1 => "11110101", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            2222 => (0 => "11110111", 1 => "11110101", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            2223 => (0 => "11110100", 1 => "11110101", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            2224 => (0 => "01110110", 1 => "11110110", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            2225 => (0 => "10110110", 1 => "11110110", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            2226 => (0 => "11010110", 1 => "11110110", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            2227 => (0 => "11100110", 1 => "11110110", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            2228 => (0 => "11111110", 1 => "11110110", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            2229 => (0 => "11110010", 1 => "11110110", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            2230 => (0 => "11110100", 1 => "11110110", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            2231 => (0 => "11110111", 1 => "11110110", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            2232 => (0 => "01110111", 1 => "11110111", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            2233 => (0 => "10110111", 1 => "11110111", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            2234 => (0 => "11010111", 1 => "11110111", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            2235 => (0 => "11100111", 1 => "11110111", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            2236 => (0 => "11111111", 1 => "11110111", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            2237 => (0 => "11110011", 1 => "11110111", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            2238 => (0 => "11110101", 1 => "11110111", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            2239 => (0 => "11110110", 1 => "11110111", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            2240 => (0 => "01111000", 1 => "11111000", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            2241 => (0 => "10111000", 1 => "11111000", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            2242 => (0 => "11011000", 1 => "11111000", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            2243 => (0 => "11101000", 1 => "11111000", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            2244 => (0 => "11110000", 1 => "11111000", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            2245 => (0 => "11111100", 1 => "11111000", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            2246 => (0 => "11111010", 1 => "11111000", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            2247 => (0 => "11111001", 1 => "11111000", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            2248 => (0 => "01111001", 1 => "11111001", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            2249 => (0 => "10111001", 1 => "11111001", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            2250 => (0 => "11011001", 1 => "11111001", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            2251 => (0 => "11101001", 1 => "11111001", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            2252 => (0 => "11110001", 1 => "11111001", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            2253 => (0 => "11111101", 1 => "11111001", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            2254 => (0 => "11111011", 1 => "11111001", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            2255 => (0 => "11111000", 1 => "11111001", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            2256 => (0 => "01111010", 1 => "11111010", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            2257 => (0 => "10111010", 1 => "11111010", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            2258 => (0 => "11011010", 1 => "11111010", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            2259 => (0 => "11101010", 1 => "11111010", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            2260 => (0 => "11110010", 1 => "11111010", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            2261 => (0 => "11111110", 1 => "11111010", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            2262 => (0 => "11111000", 1 => "11111010", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            2263 => (0 => "11111011", 1 => "11111010", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            2264 => (0 => "01111011", 1 => "11111011", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            2265 => (0 => "10111011", 1 => "11111011", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            2266 => (0 => "11011011", 1 => "11111011", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            2267 => (0 => "11101011", 1 => "11111011", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            2268 => (0 => "11110011", 1 => "11111011", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            2269 => (0 => "11111111", 1 => "11111011", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            2270 => (0 => "11111001", 1 => "11111011", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            2271 => (0 => "11111010", 1 => "11111011", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            2272 => (0 => "01111100", 1 => "11111100", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            2273 => (0 => "10111100", 1 => "11111100", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            2274 => (0 => "11011100", 1 => "11111100", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            2275 => (0 => "11101100", 1 => "11111100", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            2276 => (0 => "11110100", 1 => "11111100", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            2277 => (0 => "11111000", 1 => "11111100", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            2278 => (0 => "11111110", 1 => "11111100", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            2279 => (0 => "11111101", 1 => "11111100", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            2280 => (0 => "01111101", 1 => "11111101", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            2281 => (0 => "10111101", 1 => "11111101", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            2282 => (0 => "11011101", 1 => "11111101", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            2283 => (0 => "11101101", 1 => "11111101", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            2284 => (0 => "11110101", 1 => "11111101", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            2285 => (0 => "11111001", 1 => "11111101", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            2286 => (0 => "11111111", 1 => "11111101", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            2287 => (0 => "11111100", 1 => "11111101", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            2288 => (0 => "01111110", 1 => "11111110", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            2289 => (0 => "10111110", 1 => "11111110", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            2290 => (0 => "11011110", 1 => "11111110", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            2291 => (0 => "11101110", 1 => "11111110", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            2292 => (0 => "11110110", 1 => "11111110", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            2293 => (0 => "11111010", 1 => "11111110", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            2294 => (0 => "11111100", 1 => "11111110", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            2295 => (0 => "11111111", 1 => "11111110", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            2296 => (0 => "01111111", 1 => "11111111", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            2297 => (0 => "10111111", 1 => "11111111", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            2298 => (0 => "11011111", 1 => "11111111", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            2299 => (0 => "11101111", 1 => "11111111", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            2300 => (0 => "11110111", 1 => "11111111", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            2301 => (0 => "11111011", 1 => "11111111", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            2302 => (0 => "11111101", 1 => "11111111", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            2303 => (0 => "11111110", 1 => "11111111", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            2304 => (0 => "10000000", 1 => "01000000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            2305 => (0 => "01000000", 1 => "00100000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            2306 => (0 => "00100000", 1 => "00010000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            2307 => (0 => "00010000", 1 => "00001000", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            2308 => (0 => "00001000", 1 => "00000100", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            2309 => (0 => "00000100", 1 => "00000010", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            2310 => (0 => "00000010", 1 => "00000001", 2 => "00000000", 3 => "00000000", 4 => "11111111"),
            2311 => (0 => "10000001", 1 => "01000001", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            2312 => (0 => "01000001", 1 => "00100001", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            2313 => (0 => "00100001", 1 => "00010001", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            2314 => (0 => "00010001", 1 => "00001001", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            2315 => (0 => "00001001", 1 => "00000101", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            2316 => (0 => "00000101", 1 => "00000011", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            2317 => (0 => "00000011", 1 => "00000000", 2 => "00000001", 3 => "00000001", 4 => "11111111"),
            2318 => (0 => "10000010", 1 => "01000010", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            2319 => (0 => "01000010", 1 => "00100010", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            2320 => (0 => "00100010", 1 => "00010010", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            2321 => (0 => "00010010", 1 => "00001010", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            2322 => (0 => "00001010", 1 => "00000110", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            2323 => (0 => "00000110", 1 => "00000000", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            2324 => (0 => "00000000", 1 => "00000011", 2 => "00000010", 3 => "00000010", 4 => "11111111"),
            2325 => (0 => "10000011", 1 => "01000011", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            2326 => (0 => "01000011", 1 => "00100011", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            2327 => (0 => "00100011", 1 => "00010011", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            2328 => (0 => "00010011", 1 => "00001011", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            2329 => (0 => "00001011", 1 => "00000111", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            2330 => (0 => "00000111", 1 => "00000001", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            2331 => (0 => "00000001", 1 => "00000010", 2 => "00000011", 3 => "00000011", 4 => "11111111"),
            2332 => (0 => "10000100", 1 => "01000100", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            2333 => (0 => "01000100", 1 => "00100100", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            2334 => (0 => "00100100", 1 => "00010100", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            2335 => (0 => "00010100", 1 => "00001100", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            2336 => (0 => "00001100", 1 => "00000000", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            2337 => (0 => "00000000", 1 => "00000110", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            2338 => (0 => "00000110", 1 => "00000101", 2 => "00000100", 3 => "00000100", 4 => "11111111"),
            2339 => (0 => "10000101", 1 => "01000101", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            2340 => (0 => "01000101", 1 => "00100101", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            2341 => (0 => "00100101", 1 => "00010101", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            2342 => (0 => "00010101", 1 => "00001101", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            2343 => (0 => "00001101", 1 => "00000001", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            2344 => (0 => "00000001", 1 => "00000111", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            2345 => (0 => "00000111", 1 => "00000100", 2 => "00000101", 3 => "00000101", 4 => "11111111"),
            2346 => (0 => "10000110", 1 => "01000110", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            2347 => (0 => "01000110", 1 => "00100110", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            2348 => (0 => "00100110", 1 => "00010110", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            2349 => (0 => "00010110", 1 => "00001110", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            2350 => (0 => "00001110", 1 => "00000010", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            2351 => (0 => "00000010", 1 => "00000100", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            2352 => (0 => "00000100", 1 => "00000111", 2 => "00000110", 3 => "00000110", 4 => "11111111"),
            2353 => (0 => "10000111", 1 => "01000111", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            2354 => (0 => "01000111", 1 => "00100111", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            2355 => (0 => "00100111", 1 => "00010111", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            2356 => (0 => "00010111", 1 => "00001111", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            2357 => (0 => "00001111", 1 => "00000011", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            2358 => (0 => "00000011", 1 => "00000101", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            2359 => (0 => "00000101", 1 => "00000110", 2 => "00000111", 3 => "00000111", 4 => "11111111"),
            2360 => (0 => "10001000", 1 => "01001000", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            2361 => (0 => "01001000", 1 => "00101000", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            2362 => (0 => "00101000", 1 => "00011000", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            2363 => (0 => "00011000", 1 => "00000000", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            2364 => (0 => "00000000", 1 => "00001100", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            2365 => (0 => "00001100", 1 => "00001010", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            2366 => (0 => "00001010", 1 => "00001001", 2 => "00001000", 3 => "00001000", 4 => "11111111"),
            2367 => (0 => "10001001", 1 => "01001001", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            2368 => (0 => "01001001", 1 => "00101001", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            2369 => (0 => "00101001", 1 => "00011001", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            2370 => (0 => "00011001", 1 => "00000001", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            2371 => (0 => "00000001", 1 => "00001101", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            2372 => (0 => "00001101", 1 => "00001011", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            2373 => (0 => "00001011", 1 => "00001000", 2 => "00001001", 3 => "00001001", 4 => "11111111"),
            2374 => (0 => "10001010", 1 => "01001010", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            2375 => (0 => "01001010", 1 => "00101010", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            2376 => (0 => "00101010", 1 => "00011010", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            2377 => (0 => "00011010", 1 => "00000010", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            2378 => (0 => "00000010", 1 => "00001110", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            2379 => (0 => "00001110", 1 => "00001000", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            2380 => (0 => "00001000", 1 => "00001011", 2 => "00001010", 3 => "00001010", 4 => "11111111"),
            2381 => (0 => "10001011", 1 => "01001011", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            2382 => (0 => "01001011", 1 => "00101011", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            2383 => (0 => "00101011", 1 => "00011011", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            2384 => (0 => "00011011", 1 => "00000011", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            2385 => (0 => "00000011", 1 => "00001111", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            2386 => (0 => "00001111", 1 => "00001001", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            2387 => (0 => "00001001", 1 => "00001010", 2 => "00001011", 3 => "00001011", 4 => "11111111"),
            2388 => (0 => "10001100", 1 => "01001100", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            2389 => (0 => "01001100", 1 => "00101100", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            2390 => (0 => "00101100", 1 => "00011100", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            2391 => (0 => "00011100", 1 => "00000100", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            2392 => (0 => "00000100", 1 => "00001000", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            2393 => (0 => "00001000", 1 => "00001110", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            2394 => (0 => "00001110", 1 => "00001101", 2 => "00001100", 3 => "00001100", 4 => "11111111"),
            2395 => (0 => "10001101", 1 => "01001101", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            2396 => (0 => "01001101", 1 => "00101101", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            2397 => (0 => "00101101", 1 => "00011101", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            2398 => (0 => "00011101", 1 => "00000101", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            2399 => (0 => "00000101", 1 => "00001001", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            2400 => (0 => "00001001", 1 => "00001111", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            2401 => (0 => "00001111", 1 => "00001100", 2 => "00001101", 3 => "00001101", 4 => "11111111"),
            2402 => (0 => "10001110", 1 => "01001110", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            2403 => (0 => "01001110", 1 => "00101110", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            2404 => (0 => "00101110", 1 => "00011110", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            2405 => (0 => "00011110", 1 => "00000110", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            2406 => (0 => "00000110", 1 => "00001010", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            2407 => (0 => "00001010", 1 => "00001100", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            2408 => (0 => "00001100", 1 => "00001111", 2 => "00001110", 3 => "00001110", 4 => "11111111"),
            2409 => (0 => "10001111", 1 => "01001111", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            2410 => (0 => "01001111", 1 => "00101111", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            2411 => (0 => "00101111", 1 => "00011111", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            2412 => (0 => "00011111", 1 => "00000111", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            2413 => (0 => "00000111", 1 => "00001011", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            2414 => (0 => "00001011", 1 => "00001101", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            2415 => (0 => "00001101", 1 => "00001110", 2 => "00001111", 3 => "00001111", 4 => "11111111"),
            2416 => (0 => "10010000", 1 => "01010000", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            2417 => (0 => "01010000", 1 => "00110000", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            2418 => (0 => "00110000", 1 => "00000000", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            2419 => (0 => "00000000", 1 => "00011000", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            2420 => (0 => "00011000", 1 => "00010100", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            2421 => (0 => "00010100", 1 => "00010010", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            2422 => (0 => "00010010", 1 => "00010001", 2 => "00010000", 3 => "00010000", 4 => "11111111"),
            2423 => (0 => "10010001", 1 => "01010001", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            2424 => (0 => "01010001", 1 => "00110001", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            2425 => (0 => "00110001", 1 => "00000001", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            2426 => (0 => "00000001", 1 => "00011001", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            2427 => (0 => "00011001", 1 => "00010101", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            2428 => (0 => "00010101", 1 => "00010011", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            2429 => (0 => "00010011", 1 => "00010000", 2 => "00010001", 3 => "00010001", 4 => "11111111"),
            2430 => (0 => "10010010", 1 => "01010010", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            2431 => (0 => "01010010", 1 => "00110010", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            2432 => (0 => "00110010", 1 => "00000010", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            2433 => (0 => "00000010", 1 => "00011010", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            2434 => (0 => "00011010", 1 => "00010110", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            2435 => (0 => "00010110", 1 => "00010000", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            2436 => (0 => "00010000", 1 => "00010011", 2 => "00010010", 3 => "00010010", 4 => "11111111"),
            2437 => (0 => "10010011", 1 => "01010011", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            2438 => (0 => "01010011", 1 => "00110011", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            2439 => (0 => "00110011", 1 => "00000011", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            2440 => (0 => "00000011", 1 => "00011011", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            2441 => (0 => "00011011", 1 => "00010111", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            2442 => (0 => "00010111", 1 => "00010001", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            2443 => (0 => "00010001", 1 => "00010010", 2 => "00010011", 3 => "00010011", 4 => "11111111"),
            2444 => (0 => "10010100", 1 => "01010100", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            2445 => (0 => "01010100", 1 => "00110100", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            2446 => (0 => "00110100", 1 => "00000100", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            2447 => (0 => "00000100", 1 => "00011100", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            2448 => (0 => "00011100", 1 => "00010000", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            2449 => (0 => "00010000", 1 => "00010110", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            2450 => (0 => "00010110", 1 => "00010101", 2 => "00010100", 3 => "00010100", 4 => "11111111"),
            2451 => (0 => "10010101", 1 => "01010101", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            2452 => (0 => "01010101", 1 => "00110101", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            2453 => (0 => "00110101", 1 => "00000101", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            2454 => (0 => "00000101", 1 => "00011101", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            2455 => (0 => "00011101", 1 => "00010001", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            2456 => (0 => "00010001", 1 => "00010111", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            2457 => (0 => "00010111", 1 => "00010100", 2 => "00010101", 3 => "00010101", 4 => "11111111"),
            2458 => (0 => "10010110", 1 => "01010110", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            2459 => (0 => "01010110", 1 => "00110110", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            2460 => (0 => "00110110", 1 => "00000110", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            2461 => (0 => "00000110", 1 => "00011110", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            2462 => (0 => "00011110", 1 => "00010010", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            2463 => (0 => "00010010", 1 => "00010100", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            2464 => (0 => "00010100", 1 => "00010111", 2 => "00010110", 3 => "00010110", 4 => "11111111"),
            2465 => (0 => "10010111", 1 => "01010111", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            2466 => (0 => "01010111", 1 => "00110111", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            2467 => (0 => "00110111", 1 => "00000111", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            2468 => (0 => "00000111", 1 => "00011111", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            2469 => (0 => "00011111", 1 => "00010011", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            2470 => (0 => "00010011", 1 => "00010101", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            2471 => (0 => "00010101", 1 => "00010110", 2 => "00010111", 3 => "00010111", 4 => "11111111"),
            2472 => (0 => "10011000", 1 => "01011000", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            2473 => (0 => "01011000", 1 => "00111000", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            2474 => (0 => "00111000", 1 => "00001000", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            2475 => (0 => "00001000", 1 => "00010000", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            2476 => (0 => "00010000", 1 => "00011100", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            2477 => (0 => "00011100", 1 => "00011010", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            2478 => (0 => "00011010", 1 => "00011001", 2 => "00011000", 3 => "00011000", 4 => "11111111"),
            2479 => (0 => "10011001", 1 => "01011001", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            2480 => (0 => "01011001", 1 => "00111001", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            2481 => (0 => "00111001", 1 => "00001001", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            2482 => (0 => "00001001", 1 => "00010001", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            2483 => (0 => "00010001", 1 => "00011101", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            2484 => (0 => "00011101", 1 => "00011011", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            2485 => (0 => "00011011", 1 => "00011000", 2 => "00011001", 3 => "00011001", 4 => "11111111"),
            2486 => (0 => "10011010", 1 => "01011010", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            2487 => (0 => "01011010", 1 => "00111010", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            2488 => (0 => "00111010", 1 => "00001010", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            2489 => (0 => "00001010", 1 => "00010010", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            2490 => (0 => "00010010", 1 => "00011110", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            2491 => (0 => "00011110", 1 => "00011000", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            2492 => (0 => "00011000", 1 => "00011011", 2 => "00011010", 3 => "00011010", 4 => "11111111"),
            2493 => (0 => "10011011", 1 => "01011011", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            2494 => (0 => "01011011", 1 => "00111011", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            2495 => (0 => "00111011", 1 => "00001011", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            2496 => (0 => "00001011", 1 => "00010011", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            2497 => (0 => "00010011", 1 => "00011111", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            2498 => (0 => "00011111", 1 => "00011001", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            2499 => (0 => "00011001", 1 => "00011010", 2 => "00011011", 3 => "00011011", 4 => "11111111"),
            2500 => (0 => "10011100", 1 => "01011100", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            2501 => (0 => "01011100", 1 => "00111100", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            2502 => (0 => "00111100", 1 => "00001100", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            2503 => (0 => "00001100", 1 => "00010100", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            2504 => (0 => "00010100", 1 => "00011000", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            2505 => (0 => "00011000", 1 => "00011110", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            2506 => (0 => "00011110", 1 => "00011101", 2 => "00011100", 3 => "00011100", 4 => "11111111"),
            2507 => (0 => "10011101", 1 => "01011101", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            2508 => (0 => "01011101", 1 => "00111101", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            2509 => (0 => "00111101", 1 => "00001101", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            2510 => (0 => "00001101", 1 => "00010101", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            2511 => (0 => "00010101", 1 => "00011001", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            2512 => (0 => "00011001", 1 => "00011111", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            2513 => (0 => "00011111", 1 => "00011100", 2 => "00011101", 3 => "00011101", 4 => "11111111"),
            2514 => (0 => "10011110", 1 => "01011110", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            2515 => (0 => "01011110", 1 => "00111110", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            2516 => (0 => "00111110", 1 => "00001110", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            2517 => (0 => "00001110", 1 => "00010110", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            2518 => (0 => "00010110", 1 => "00011010", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            2519 => (0 => "00011010", 1 => "00011100", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            2520 => (0 => "00011100", 1 => "00011111", 2 => "00011110", 3 => "00011110", 4 => "11111111"),
            2521 => (0 => "10011111", 1 => "01011111", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            2522 => (0 => "01011111", 1 => "00111111", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            2523 => (0 => "00111111", 1 => "00001111", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            2524 => (0 => "00001111", 1 => "00010111", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            2525 => (0 => "00010111", 1 => "00011011", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            2526 => (0 => "00011011", 1 => "00011101", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            2527 => (0 => "00011101", 1 => "00011110", 2 => "00011111", 3 => "00011111", 4 => "11111111"),
            2528 => (0 => "10100000", 1 => "01100000", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            2529 => (0 => "01100000", 1 => "00000000", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            2530 => (0 => "00000000", 1 => "00110000", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            2531 => (0 => "00110000", 1 => "00101000", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            2532 => (0 => "00101000", 1 => "00100100", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            2533 => (0 => "00100100", 1 => "00100010", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            2534 => (0 => "00100010", 1 => "00100001", 2 => "00100000", 3 => "00100000", 4 => "11111111"),
            2535 => (0 => "10100001", 1 => "01100001", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            2536 => (0 => "01100001", 1 => "00000001", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            2537 => (0 => "00000001", 1 => "00110001", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            2538 => (0 => "00110001", 1 => "00101001", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            2539 => (0 => "00101001", 1 => "00100101", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            2540 => (0 => "00100101", 1 => "00100011", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            2541 => (0 => "00100011", 1 => "00100000", 2 => "00100001", 3 => "00100001", 4 => "11111111"),
            2542 => (0 => "10100010", 1 => "01100010", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            2543 => (0 => "01100010", 1 => "00000010", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            2544 => (0 => "00000010", 1 => "00110010", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            2545 => (0 => "00110010", 1 => "00101010", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            2546 => (0 => "00101010", 1 => "00100110", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            2547 => (0 => "00100110", 1 => "00100000", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            2548 => (0 => "00100000", 1 => "00100011", 2 => "00100010", 3 => "00100010", 4 => "11111111"),
            2549 => (0 => "10100011", 1 => "01100011", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            2550 => (0 => "01100011", 1 => "00000011", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            2551 => (0 => "00000011", 1 => "00110011", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            2552 => (0 => "00110011", 1 => "00101011", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            2553 => (0 => "00101011", 1 => "00100111", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            2554 => (0 => "00100111", 1 => "00100001", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            2555 => (0 => "00100001", 1 => "00100010", 2 => "00100011", 3 => "00100011", 4 => "11111111"),
            2556 => (0 => "10100100", 1 => "01100100", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            2557 => (0 => "01100100", 1 => "00000100", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            2558 => (0 => "00000100", 1 => "00110100", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            2559 => (0 => "00110100", 1 => "00101100", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            2560 => (0 => "00101100", 1 => "00100000", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            2561 => (0 => "00100000", 1 => "00100110", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            2562 => (0 => "00100110", 1 => "00100101", 2 => "00100100", 3 => "00100100", 4 => "11111111"),
            2563 => (0 => "10100101", 1 => "01100101", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            2564 => (0 => "01100101", 1 => "00000101", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            2565 => (0 => "00000101", 1 => "00110101", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            2566 => (0 => "00110101", 1 => "00101101", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            2567 => (0 => "00101101", 1 => "00100001", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            2568 => (0 => "00100001", 1 => "00100111", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            2569 => (0 => "00100111", 1 => "00100100", 2 => "00100101", 3 => "00100101", 4 => "11111111"),
            2570 => (0 => "10100110", 1 => "01100110", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            2571 => (0 => "01100110", 1 => "00000110", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            2572 => (0 => "00000110", 1 => "00110110", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            2573 => (0 => "00110110", 1 => "00101110", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            2574 => (0 => "00101110", 1 => "00100010", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            2575 => (0 => "00100010", 1 => "00100100", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            2576 => (0 => "00100100", 1 => "00100111", 2 => "00100110", 3 => "00100110", 4 => "11111111"),
            2577 => (0 => "10100111", 1 => "01100111", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            2578 => (0 => "01100111", 1 => "00000111", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            2579 => (0 => "00000111", 1 => "00110111", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            2580 => (0 => "00110111", 1 => "00101111", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            2581 => (0 => "00101111", 1 => "00100011", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            2582 => (0 => "00100011", 1 => "00100101", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            2583 => (0 => "00100101", 1 => "00100110", 2 => "00100111", 3 => "00100111", 4 => "11111111"),
            2584 => (0 => "10101000", 1 => "01101000", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            2585 => (0 => "01101000", 1 => "00001000", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            2586 => (0 => "00001000", 1 => "00111000", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            2587 => (0 => "00111000", 1 => "00100000", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            2588 => (0 => "00100000", 1 => "00101100", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            2589 => (0 => "00101100", 1 => "00101010", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            2590 => (0 => "00101010", 1 => "00101001", 2 => "00101000", 3 => "00101000", 4 => "11111111"),
            2591 => (0 => "10101001", 1 => "01101001", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            2592 => (0 => "01101001", 1 => "00001001", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            2593 => (0 => "00001001", 1 => "00111001", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            2594 => (0 => "00111001", 1 => "00100001", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            2595 => (0 => "00100001", 1 => "00101101", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            2596 => (0 => "00101101", 1 => "00101011", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            2597 => (0 => "00101011", 1 => "00101000", 2 => "00101001", 3 => "00101001", 4 => "11111111"),
            2598 => (0 => "10101010", 1 => "01101010", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            2599 => (0 => "01101010", 1 => "00001010", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            2600 => (0 => "00001010", 1 => "00111010", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            2601 => (0 => "00111010", 1 => "00100010", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            2602 => (0 => "00100010", 1 => "00101110", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            2603 => (0 => "00101110", 1 => "00101000", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            2604 => (0 => "00101000", 1 => "00101011", 2 => "00101010", 3 => "00101010", 4 => "11111111"),
            2605 => (0 => "10101011", 1 => "01101011", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            2606 => (0 => "01101011", 1 => "00001011", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            2607 => (0 => "00001011", 1 => "00111011", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            2608 => (0 => "00111011", 1 => "00100011", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            2609 => (0 => "00100011", 1 => "00101111", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            2610 => (0 => "00101111", 1 => "00101001", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            2611 => (0 => "00101001", 1 => "00101010", 2 => "00101011", 3 => "00101011", 4 => "11111111"),
            2612 => (0 => "10101100", 1 => "01101100", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            2613 => (0 => "01101100", 1 => "00001100", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            2614 => (0 => "00001100", 1 => "00111100", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            2615 => (0 => "00111100", 1 => "00100100", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            2616 => (0 => "00100100", 1 => "00101000", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            2617 => (0 => "00101000", 1 => "00101110", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            2618 => (0 => "00101110", 1 => "00101101", 2 => "00101100", 3 => "00101100", 4 => "11111111"),
            2619 => (0 => "10101101", 1 => "01101101", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            2620 => (0 => "01101101", 1 => "00001101", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            2621 => (0 => "00001101", 1 => "00111101", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            2622 => (0 => "00111101", 1 => "00100101", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            2623 => (0 => "00100101", 1 => "00101001", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            2624 => (0 => "00101001", 1 => "00101111", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            2625 => (0 => "00101111", 1 => "00101100", 2 => "00101101", 3 => "00101101", 4 => "11111111"),
            2626 => (0 => "10101110", 1 => "01101110", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            2627 => (0 => "01101110", 1 => "00001110", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            2628 => (0 => "00001110", 1 => "00111110", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            2629 => (0 => "00111110", 1 => "00100110", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            2630 => (0 => "00100110", 1 => "00101010", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            2631 => (0 => "00101010", 1 => "00101100", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            2632 => (0 => "00101100", 1 => "00101111", 2 => "00101110", 3 => "00101110", 4 => "11111111"),
            2633 => (0 => "10101111", 1 => "01101111", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            2634 => (0 => "01101111", 1 => "00001111", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            2635 => (0 => "00001111", 1 => "00111111", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            2636 => (0 => "00111111", 1 => "00100111", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            2637 => (0 => "00100111", 1 => "00101011", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            2638 => (0 => "00101011", 1 => "00101101", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            2639 => (0 => "00101101", 1 => "00101110", 2 => "00101111", 3 => "00101111", 4 => "11111111"),
            2640 => (0 => "10110000", 1 => "01110000", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            2641 => (0 => "01110000", 1 => "00010000", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            2642 => (0 => "00010000", 1 => "00100000", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            2643 => (0 => "00100000", 1 => "00111000", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            2644 => (0 => "00111000", 1 => "00110100", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            2645 => (0 => "00110100", 1 => "00110010", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            2646 => (0 => "00110010", 1 => "00110001", 2 => "00110000", 3 => "00110000", 4 => "11111111"),
            2647 => (0 => "10110001", 1 => "01110001", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            2648 => (0 => "01110001", 1 => "00010001", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            2649 => (0 => "00010001", 1 => "00100001", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            2650 => (0 => "00100001", 1 => "00111001", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            2651 => (0 => "00111001", 1 => "00110101", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            2652 => (0 => "00110101", 1 => "00110011", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            2653 => (0 => "00110011", 1 => "00110000", 2 => "00110001", 3 => "00110001", 4 => "11111111"),
            2654 => (0 => "10110010", 1 => "01110010", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            2655 => (0 => "01110010", 1 => "00010010", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            2656 => (0 => "00010010", 1 => "00100010", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            2657 => (0 => "00100010", 1 => "00111010", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            2658 => (0 => "00111010", 1 => "00110110", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            2659 => (0 => "00110110", 1 => "00110000", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            2660 => (0 => "00110000", 1 => "00110011", 2 => "00110010", 3 => "00110010", 4 => "11111111"),
            2661 => (0 => "10110011", 1 => "01110011", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            2662 => (0 => "01110011", 1 => "00010011", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            2663 => (0 => "00010011", 1 => "00100011", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            2664 => (0 => "00100011", 1 => "00111011", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            2665 => (0 => "00111011", 1 => "00110111", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            2666 => (0 => "00110111", 1 => "00110001", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            2667 => (0 => "00110001", 1 => "00110010", 2 => "00110011", 3 => "00110011", 4 => "11111111"),
            2668 => (0 => "10110100", 1 => "01110100", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            2669 => (0 => "01110100", 1 => "00010100", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            2670 => (0 => "00010100", 1 => "00100100", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            2671 => (0 => "00100100", 1 => "00111100", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            2672 => (0 => "00111100", 1 => "00110000", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            2673 => (0 => "00110000", 1 => "00110110", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            2674 => (0 => "00110110", 1 => "00110101", 2 => "00110100", 3 => "00110100", 4 => "11111111"),
            2675 => (0 => "10110101", 1 => "01110101", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            2676 => (0 => "01110101", 1 => "00010101", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            2677 => (0 => "00010101", 1 => "00100101", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            2678 => (0 => "00100101", 1 => "00111101", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            2679 => (0 => "00111101", 1 => "00110001", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            2680 => (0 => "00110001", 1 => "00110111", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            2681 => (0 => "00110111", 1 => "00110100", 2 => "00110101", 3 => "00110101", 4 => "11111111"),
            2682 => (0 => "10110110", 1 => "01110110", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            2683 => (0 => "01110110", 1 => "00010110", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            2684 => (0 => "00010110", 1 => "00100110", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            2685 => (0 => "00100110", 1 => "00111110", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            2686 => (0 => "00111110", 1 => "00110010", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            2687 => (0 => "00110010", 1 => "00110100", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            2688 => (0 => "00110100", 1 => "00110111", 2 => "00110110", 3 => "00110110", 4 => "11111111"),
            2689 => (0 => "10110111", 1 => "01110111", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            2690 => (0 => "01110111", 1 => "00010111", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            2691 => (0 => "00010111", 1 => "00100111", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            2692 => (0 => "00100111", 1 => "00111111", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            2693 => (0 => "00111111", 1 => "00110011", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            2694 => (0 => "00110011", 1 => "00110101", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            2695 => (0 => "00110101", 1 => "00110110", 2 => "00110111", 3 => "00110111", 4 => "11111111"),
            2696 => (0 => "10111000", 1 => "01111000", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            2697 => (0 => "01111000", 1 => "00011000", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            2698 => (0 => "00011000", 1 => "00101000", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            2699 => (0 => "00101000", 1 => "00110000", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            2700 => (0 => "00110000", 1 => "00111100", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            2701 => (0 => "00111100", 1 => "00111010", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            2702 => (0 => "00111010", 1 => "00111001", 2 => "00111000", 3 => "00111000", 4 => "11111111"),
            2703 => (0 => "10111001", 1 => "01111001", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            2704 => (0 => "01111001", 1 => "00011001", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            2705 => (0 => "00011001", 1 => "00101001", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            2706 => (0 => "00101001", 1 => "00110001", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            2707 => (0 => "00110001", 1 => "00111101", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            2708 => (0 => "00111101", 1 => "00111011", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            2709 => (0 => "00111011", 1 => "00111000", 2 => "00111001", 3 => "00111001", 4 => "11111111"),
            2710 => (0 => "10111010", 1 => "01111010", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            2711 => (0 => "01111010", 1 => "00011010", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            2712 => (0 => "00011010", 1 => "00101010", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            2713 => (0 => "00101010", 1 => "00110010", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            2714 => (0 => "00110010", 1 => "00111110", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            2715 => (0 => "00111110", 1 => "00111000", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            2716 => (0 => "00111000", 1 => "00111011", 2 => "00111010", 3 => "00111010", 4 => "11111111"),
            2717 => (0 => "10111011", 1 => "01111011", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            2718 => (0 => "01111011", 1 => "00011011", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            2719 => (0 => "00011011", 1 => "00101011", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            2720 => (0 => "00101011", 1 => "00110011", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            2721 => (0 => "00110011", 1 => "00111111", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            2722 => (0 => "00111111", 1 => "00111001", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            2723 => (0 => "00111001", 1 => "00111010", 2 => "00111011", 3 => "00111011", 4 => "11111111"),
            2724 => (0 => "10111100", 1 => "01111100", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            2725 => (0 => "01111100", 1 => "00011100", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            2726 => (0 => "00011100", 1 => "00101100", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            2727 => (0 => "00101100", 1 => "00110100", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            2728 => (0 => "00110100", 1 => "00111000", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            2729 => (0 => "00111000", 1 => "00111110", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            2730 => (0 => "00111110", 1 => "00111101", 2 => "00111100", 3 => "00111100", 4 => "11111111"),
            2731 => (0 => "10111101", 1 => "01111101", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            2732 => (0 => "01111101", 1 => "00011101", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            2733 => (0 => "00011101", 1 => "00101101", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            2734 => (0 => "00101101", 1 => "00110101", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            2735 => (0 => "00110101", 1 => "00111001", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            2736 => (0 => "00111001", 1 => "00111111", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            2737 => (0 => "00111111", 1 => "00111100", 2 => "00111101", 3 => "00111101", 4 => "11111111"),
            2738 => (0 => "10111110", 1 => "01111110", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            2739 => (0 => "01111110", 1 => "00011110", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            2740 => (0 => "00011110", 1 => "00101110", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            2741 => (0 => "00101110", 1 => "00110110", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            2742 => (0 => "00110110", 1 => "00111010", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            2743 => (0 => "00111010", 1 => "00111100", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            2744 => (0 => "00111100", 1 => "00111111", 2 => "00111110", 3 => "00111110", 4 => "11111111"),
            2745 => (0 => "10111111", 1 => "01111111", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            2746 => (0 => "01111111", 1 => "00011111", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            2747 => (0 => "00011111", 1 => "00101111", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            2748 => (0 => "00101111", 1 => "00110111", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            2749 => (0 => "00110111", 1 => "00111011", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            2750 => (0 => "00111011", 1 => "00111101", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            2751 => (0 => "00111101", 1 => "00111110", 2 => "00111111", 3 => "00111111", 4 => "11111111"),
            2752 => (0 => "11000000", 1 => "00000000", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            2753 => (0 => "00000000", 1 => "01100000", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            2754 => (0 => "01100000", 1 => "01010000", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            2755 => (0 => "01010000", 1 => "01001000", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            2756 => (0 => "01001000", 1 => "01000100", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            2757 => (0 => "01000100", 1 => "01000010", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            2758 => (0 => "01000010", 1 => "01000001", 2 => "01000000", 3 => "01000000", 4 => "11111111"),
            2759 => (0 => "11000001", 1 => "00000001", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            2760 => (0 => "00000001", 1 => "01100001", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            2761 => (0 => "01100001", 1 => "01010001", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            2762 => (0 => "01010001", 1 => "01001001", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            2763 => (0 => "01001001", 1 => "01000101", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            2764 => (0 => "01000101", 1 => "01000011", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            2765 => (0 => "01000011", 1 => "01000000", 2 => "01000001", 3 => "01000001", 4 => "11111111"),
            2766 => (0 => "11000010", 1 => "00000010", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            2767 => (0 => "00000010", 1 => "01100010", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            2768 => (0 => "01100010", 1 => "01010010", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            2769 => (0 => "01010010", 1 => "01001010", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            2770 => (0 => "01001010", 1 => "01000110", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            2771 => (0 => "01000110", 1 => "01000000", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            2772 => (0 => "01000000", 1 => "01000011", 2 => "01000010", 3 => "01000010", 4 => "11111111"),
            2773 => (0 => "11000011", 1 => "00000011", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            2774 => (0 => "00000011", 1 => "01100011", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            2775 => (0 => "01100011", 1 => "01010011", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            2776 => (0 => "01010011", 1 => "01001011", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            2777 => (0 => "01001011", 1 => "01000111", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            2778 => (0 => "01000111", 1 => "01000001", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            2779 => (0 => "01000001", 1 => "01000010", 2 => "01000011", 3 => "01000011", 4 => "11111111"),
            2780 => (0 => "11000100", 1 => "00000100", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            2781 => (0 => "00000100", 1 => "01100100", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            2782 => (0 => "01100100", 1 => "01010100", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            2783 => (0 => "01010100", 1 => "01001100", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            2784 => (0 => "01001100", 1 => "01000000", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            2785 => (0 => "01000000", 1 => "01000110", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            2786 => (0 => "01000110", 1 => "01000101", 2 => "01000100", 3 => "01000100", 4 => "11111111"),
            2787 => (0 => "11000101", 1 => "00000101", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            2788 => (0 => "00000101", 1 => "01100101", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            2789 => (0 => "01100101", 1 => "01010101", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            2790 => (0 => "01010101", 1 => "01001101", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            2791 => (0 => "01001101", 1 => "01000001", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            2792 => (0 => "01000001", 1 => "01000111", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            2793 => (0 => "01000111", 1 => "01000100", 2 => "01000101", 3 => "01000101", 4 => "11111111"),
            2794 => (0 => "11000110", 1 => "00000110", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            2795 => (0 => "00000110", 1 => "01100110", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            2796 => (0 => "01100110", 1 => "01010110", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            2797 => (0 => "01010110", 1 => "01001110", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            2798 => (0 => "01001110", 1 => "01000010", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            2799 => (0 => "01000010", 1 => "01000100", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            2800 => (0 => "01000100", 1 => "01000111", 2 => "01000110", 3 => "01000110", 4 => "11111111"),
            2801 => (0 => "11000111", 1 => "00000111", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            2802 => (0 => "00000111", 1 => "01100111", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            2803 => (0 => "01100111", 1 => "01010111", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            2804 => (0 => "01010111", 1 => "01001111", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            2805 => (0 => "01001111", 1 => "01000011", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            2806 => (0 => "01000011", 1 => "01000101", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            2807 => (0 => "01000101", 1 => "01000110", 2 => "01000111", 3 => "01000111", 4 => "11111111"),
            2808 => (0 => "11001000", 1 => "00001000", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            2809 => (0 => "00001000", 1 => "01101000", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            2810 => (0 => "01101000", 1 => "01011000", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            2811 => (0 => "01011000", 1 => "01000000", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            2812 => (0 => "01000000", 1 => "01001100", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            2813 => (0 => "01001100", 1 => "01001010", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            2814 => (0 => "01001010", 1 => "01001001", 2 => "01001000", 3 => "01001000", 4 => "11111111"),
            2815 => (0 => "11001001", 1 => "00001001", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            2816 => (0 => "00001001", 1 => "01101001", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            2817 => (0 => "01101001", 1 => "01011001", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            2818 => (0 => "01011001", 1 => "01000001", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            2819 => (0 => "01000001", 1 => "01001101", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            2820 => (0 => "01001101", 1 => "01001011", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            2821 => (0 => "01001011", 1 => "01001000", 2 => "01001001", 3 => "01001001", 4 => "11111111"),
            2822 => (0 => "11001010", 1 => "00001010", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            2823 => (0 => "00001010", 1 => "01101010", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            2824 => (0 => "01101010", 1 => "01011010", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            2825 => (0 => "01011010", 1 => "01000010", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            2826 => (0 => "01000010", 1 => "01001110", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            2827 => (0 => "01001110", 1 => "01001000", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            2828 => (0 => "01001000", 1 => "01001011", 2 => "01001010", 3 => "01001010", 4 => "11111111"),
            2829 => (0 => "11001011", 1 => "00001011", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            2830 => (0 => "00001011", 1 => "01101011", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            2831 => (0 => "01101011", 1 => "01011011", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            2832 => (0 => "01011011", 1 => "01000011", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            2833 => (0 => "01000011", 1 => "01001111", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            2834 => (0 => "01001111", 1 => "01001001", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            2835 => (0 => "01001001", 1 => "01001010", 2 => "01001011", 3 => "01001011", 4 => "11111111"),
            2836 => (0 => "11001100", 1 => "00001100", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            2837 => (0 => "00001100", 1 => "01101100", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            2838 => (0 => "01101100", 1 => "01011100", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            2839 => (0 => "01011100", 1 => "01000100", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            2840 => (0 => "01000100", 1 => "01001000", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            2841 => (0 => "01001000", 1 => "01001110", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            2842 => (0 => "01001110", 1 => "01001101", 2 => "01001100", 3 => "01001100", 4 => "11111111"),
            2843 => (0 => "11001101", 1 => "00001101", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            2844 => (0 => "00001101", 1 => "01101101", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            2845 => (0 => "01101101", 1 => "01011101", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            2846 => (0 => "01011101", 1 => "01000101", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            2847 => (0 => "01000101", 1 => "01001001", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            2848 => (0 => "01001001", 1 => "01001111", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            2849 => (0 => "01001111", 1 => "01001100", 2 => "01001101", 3 => "01001101", 4 => "11111111"),
            2850 => (0 => "11001110", 1 => "00001110", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            2851 => (0 => "00001110", 1 => "01101110", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            2852 => (0 => "01101110", 1 => "01011110", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            2853 => (0 => "01011110", 1 => "01000110", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            2854 => (0 => "01000110", 1 => "01001010", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            2855 => (0 => "01001010", 1 => "01001100", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            2856 => (0 => "01001100", 1 => "01001111", 2 => "01001110", 3 => "01001110", 4 => "11111111"),
            2857 => (0 => "11001111", 1 => "00001111", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            2858 => (0 => "00001111", 1 => "01101111", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            2859 => (0 => "01101111", 1 => "01011111", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            2860 => (0 => "01011111", 1 => "01000111", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            2861 => (0 => "01000111", 1 => "01001011", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            2862 => (0 => "01001011", 1 => "01001101", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            2863 => (0 => "01001101", 1 => "01001110", 2 => "01001111", 3 => "01001111", 4 => "11111111"),
            2864 => (0 => "11010000", 1 => "00010000", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            2865 => (0 => "00010000", 1 => "01110000", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            2866 => (0 => "01110000", 1 => "01000000", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            2867 => (0 => "01000000", 1 => "01011000", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            2868 => (0 => "01011000", 1 => "01010100", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            2869 => (0 => "01010100", 1 => "01010010", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            2870 => (0 => "01010010", 1 => "01010001", 2 => "01010000", 3 => "01010000", 4 => "11111111"),
            2871 => (0 => "11010001", 1 => "00010001", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            2872 => (0 => "00010001", 1 => "01110001", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            2873 => (0 => "01110001", 1 => "01000001", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            2874 => (0 => "01000001", 1 => "01011001", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            2875 => (0 => "01011001", 1 => "01010101", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            2876 => (0 => "01010101", 1 => "01010011", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            2877 => (0 => "01010011", 1 => "01010000", 2 => "01010001", 3 => "01010001", 4 => "11111111"),
            2878 => (0 => "11010010", 1 => "00010010", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            2879 => (0 => "00010010", 1 => "01110010", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            2880 => (0 => "01110010", 1 => "01000010", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            2881 => (0 => "01000010", 1 => "01011010", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            2882 => (0 => "01011010", 1 => "01010110", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            2883 => (0 => "01010110", 1 => "01010000", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            2884 => (0 => "01010000", 1 => "01010011", 2 => "01010010", 3 => "01010010", 4 => "11111111"),
            2885 => (0 => "11010011", 1 => "00010011", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            2886 => (0 => "00010011", 1 => "01110011", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            2887 => (0 => "01110011", 1 => "01000011", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            2888 => (0 => "01000011", 1 => "01011011", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            2889 => (0 => "01011011", 1 => "01010111", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            2890 => (0 => "01010111", 1 => "01010001", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            2891 => (0 => "01010001", 1 => "01010010", 2 => "01010011", 3 => "01010011", 4 => "11111111"),
            2892 => (0 => "11010100", 1 => "00010100", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            2893 => (0 => "00010100", 1 => "01110100", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            2894 => (0 => "01110100", 1 => "01000100", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            2895 => (0 => "01000100", 1 => "01011100", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            2896 => (0 => "01011100", 1 => "01010000", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            2897 => (0 => "01010000", 1 => "01010110", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            2898 => (0 => "01010110", 1 => "01010101", 2 => "01010100", 3 => "01010100", 4 => "11111111"),
            2899 => (0 => "11010101", 1 => "00010101", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            2900 => (0 => "00010101", 1 => "01110101", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            2901 => (0 => "01110101", 1 => "01000101", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            2902 => (0 => "01000101", 1 => "01011101", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            2903 => (0 => "01011101", 1 => "01010001", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            2904 => (0 => "01010001", 1 => "01010111", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            2905 => (0 => "01010111", 1 => "01010100", 2 => "01010101", 3 => "01010101", 4 => "11111111"),
            2906 => (0 => "11010110", 1 => "00010110", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            2907 => (0 => "00010110", 1 => "01110110", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            2908 => (0 => "01110110", 1 => "01000110", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            2909 => (0 => "01000110", 1 => "01011110", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            2910 => (0 => "01011110", 1 => "01010010", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            2911 => (0 => "01010010", 1 => "01010100", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            2912 => (0 => "01010100", 1 => "01010111", 2 => "01010110", 3 => "01010110", 4 => "11111111"),
            2913 => (0 => "11010111", 1 => "00010111", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            2914 => (0 => "00010111", 1 => "01110111", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            2915 => (0 => "01110111", 1 => "01000111", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            2916 => (0 => "01000111", 1 => "01011111", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            2917 => (0 => "01011111", 1 => "01010011", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            2918 => (0 => "01010011", 1 => "01010101", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            2919 => (0 => "01010101", 1 => "01010110", 2 => "01010111", 3 => "01010111", 4 => "11111111"),
            2920 => (0 => "11011000", 1 => "00011000", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            2921 => (0 => "00011000", 1 => "01111000", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            2922 => (0 => "01111000", 1 => "01001000", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            2923 => (0 => "01001000", 1 => "01010000", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            2924 => (0 => "01010000", 1 => "01011100", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            2925 => (0 => "01011100", 1 => "01011010", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            2926 => (0 => "01011010", 1 => "01011001", 2 => "01011000", 3 => "01011000", 4 => "11111111"),
            2927 => (0 => "11011001", 1 => "00011001", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            2928 => (0 => "00011001", 1 => "01111001", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            2929 => (0 => "01111001", 1 => "01001001", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            2930 => (0 => "01001001", 1 => "01010001", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            2931 => (0 => "01010001", 1 => "01011101", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            2932 => (0 => "01011101", 1 => "01011011", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            2933 => (0 => "01011011", 1 => "01011000", 2 => "01011001", 3 => "01011001", 4 => "11111111"),
            2934 => (0 => "11011010", 1 => "00011010", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            2935 => (0 => "00011010", 1 => "01111010", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            2936 => (0 => "01111010", 1 => "01001010", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            2937 => (0 => "01001010", 1 => "01010010", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            2938 => (0 => "01010010", 1 => "01011110", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            2939 => (0 => "01011110", 1 => "01011000", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            2940 => (0 => "01011000", 1 => "01011011", 2 => "01011010", 3 => "01011010", 4 => "11111111"),
            2941 => (0 => "11011011", 1 => "00011011", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            2942 => (0 => "00011011", 1 => "01111011", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            2943 => (0 => "01111011", 1 => "01001011", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            2944 => (0 => "01001011", 1 => "01010011", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            2945 => (0 => "01010011", 1 => "01011111", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            2946 => (0 => "01011111", 1 => "01011001", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            2947 => (0 => "01011001", 1 => "01011010", 2 => "01011011", 3 => "01011011", 4 => "11111111"),
            2948 => (0 => "11011100", 1 => "00011100", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            2949 => (0 => "00011100", 1 => "01111100", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            2950 => (0 => "01111100", 1 => "01001100", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            2951 => (0 => "01001100", 1 => "01010100", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            2952 => (0 => "01010100", 1 => "01011000", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            2953 => (0 => "01011000", 1 => "01011110", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            2954 => (0 => "01011110", 1 => "01011101", 2 => "01011100", 3 => "01011100", 4 => "11111111"),
            2955 => (0 => "11011101", 1 => "00011101", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            2956 => (0 => "00011101", 1 => "01111101", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            2957 => (0 => "01111101", 1 => "01001101", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            2958 => (0 => "01001101", 1 => "01010101", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            2959 => (0 => "01010101", 1 => "01011001", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            2960 => (0 => "01011001", 1 => "01011111", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            2961 => (0 => "01011111", 1 => "01011100", 2 => "01011101", 3 => "01011101", 4 => "11111111"),
            2962 => (0 => "11011110", 1 => "00011110", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            2963 => (0 => "00011110", 1 => "01111110", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            2964 => (0 => "01111110", 1 => "01001110", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            2965 => (0 => "01001110", 1 => "01010110", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            2966 => (0 => "01010110", 1 => "01011010", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            2967 => (0 => "01011010", 1 => "01011100", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            2968 => (0 => "01011100", 1 => "01011111", 2 => "01011110", 3 => "01011110", 4 => "11111111"),
            2969 => (0 => "11011111", 1 => "00011111", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            2970 => (0 => "00011111", 1 => "01111111", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            2971 => (0 => "01111111", 1 => "01001111", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            2972 => (0 => "01001111", 1 => "01010111", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            2973 => (0 => "01010111", 1 => "01011011", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            2974 => (0 => "01011011", 1 => "01011101", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            2975 => (0 => "01011101", 1 => "01011110", 2 => "01011111", 3 => "01011111", 4 => "11111111"),
            2976 => (0 => "11100000", 1 => "00100000", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            2977 => (0 => "00100000", 1 => "01000000", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            2978 => (0 => "01000000", 1 => "01110000", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            2979 => (0 => "01110000", 1 => "01101000", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            2980 => (0 => "01101000", 1 => "01100100", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            2981 => (0 => "01100100", 1 => "01100010", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            2982 => (0 => "01100010", 1 => "01100001", 2 => "01100000", 3 => "01100000", 4 => "11111111"),
            2983 => (0 => "11100001", 1 => "00100001", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            2984 => (0 => "00100001", 1 => "01000001", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            2985 => (0 => "01000001", 1 => "01110001", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            2986 => (0 => "01110001", 1 => "01101001", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            2987 => (0 => "01101001", 1 => "01100101", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            2988 => (0 => "01100101", 1 => "01100011", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            2989 => (0 => "01100011", 1 => "01100000", 2 => "01100001", 3 => "01100001", 4 => "11111111"),
            2990 => (0 => "11100010", 1 => "00100010", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            2991 => (0 => "00100010", 1 => "01000010", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            2992 => (0 => "01000010", 1 => "01110010", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            2993 => (0 => "01110010", 1 => "01101010", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            2994 => (0 => "01101010", 1 => "01100110", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            2995 => (0 => "01100110", 1 => "01100000", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            2996 => (0 => "01100000", 1 => "01100011", 2 => "01100010", 3 => "01100010", 4 => "11111111"),
            2997 => (0 => "11100011", 1 => "00100011", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            2998 => (0 => "00100011", 1 => "01000011", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            2999 => (0 => "01000011", 1 => "01110011", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            3000 => (0 => "01110011", 1 => "01101011", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            3001 => (0 => "01101011", 1 => "01100111", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            3002 => (0 => "01100111", 1 => "01100001", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            3003 => (0 => "01100001", 1 => "01100010", 2 => "01100011", 3 => "01100011", 4 => "11111111"),
            3004 => (0 => "11100100", 1 => "00100100", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            3005 => (0 => "00100100", 1 => "01000100", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            3006 => (0 => "01000100", 1 => "01110100", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            3007 => (0 => "01110100", 1 => "01101100", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            3008 => (0 => "01101100", 1 => "01100000", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            3009 => (0 => "01100000", 1 => "01100110", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            3010 => (0 => "01100110", 1 => "01100101", 2 => "01100100", 3 => "01100100", 4 => "11111111"),
            3011 => (0 => "11100101", 1 => "00100101", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            3012 => (0 => "00100101", 1 => "01000101", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            3013 => (0 => "01000101", 1 => "01110101", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            3014 => (0 => "01110101", 1 => "01101101", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            3015 => (0 => "01101101", 1 => "01100001", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            3016 => (0 => "01100001", 1 => "01100111", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            3017 => (0 => "01100111", 1 => "01100100", 2 => "01100101", 3 => "01100101", 4 => "11111111"),
            3018 => (0 => "11100110", 1 => "00100110", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            3019 => (0 => "00100110", 1 => "01000110", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            3020 => (0 => "01000110", 1 => "01110110", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            3021 => (0 => "01110110", 1 => "01101110", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            3022 => (0 => "01101110", 1 => "01100010", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            3023 => (0 => "01100010", 1 => "01100100", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            3024 => (0 => "01100100", 1 => "01100111", 2 => "01100110", 3 => "01100110", 4 => "11111111"),
            3025 => (0 => "11100111", 1 => "00100111", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            3026 => (0 => "00100111", 1 => "01000111", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            3027 => (0 => "01000111", 1 => "01110111", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            3028 => (0 => "01110111", 1 => "01101111", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            3029 => (0 => "01101111", 1 => "01100011", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            3030 => (0 => "01100011", 1 => "01100101", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            3031 => (0 => "01100101", 1 => "01100110", 2 => "01100111", 3 => "01100111", 4 => "11111111"),
            3032 => (0 => "11101000", 1 => "00101000", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            3033 => (0 => "00101000", 1 => "01001000", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            3034 => (0 => "01001000", 1 => "01111000", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            3035 => (0 => "01111000", 1 => "01100000", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            3036 => (0 => "01100000", 1 => "01101100", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            3037 => (0 => "01101100", 1 => "01101010", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            3038 => (0 => "01101010", 1 => "01101001", 2 => "01101000", 3 => "01101000", 4 => "11111111"),
            3039 => (0 => "11101001", 1 => "00101001", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            3040 => (0 => "00101001", 1 => "01001001", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            3041 => (0 => "01001001", 1 => "01111001", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            3042 => (0 => "01111001", 1 => "01100001", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            3043 => (0 => "01100001", 1 => "01101101", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            3044 => (0 => "01101101", 1 => "01101011", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            3045 => (0 => "01101011", 1 => "01101000", 2 => "01101001", 3 => "01101001", 4 => "11111111"),
            3046 => (0 => "11101010", 1 => "00101010", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            3047 => (0 => "00101010", 1 => "01001010", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            3048 => (0 => "01001010", 1 => "01111010", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            3049 => (0 => "01111010", 1 => "01100010", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            3050 => (0 => "01100010", 1 => "01101110", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            3051 => (0 => "01101110", 1 => "01101000", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            3052 => (0 => "01101000", 1 => "01101011", 2 => "01101010", 3 => "01101010", 4 => "11111111"),
            3053 => (0 => "11101011", 1 => "00101011", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            3054 => (0 => "00101011", 1 => "01001011", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            3055 => (0 => "01001011", 1 => "01111011", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            3056 => (0 => "01111011", 1 => "01100011", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            3057 => (0 => "01100011", 1 => "01101111", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            3058 => (0 => "01101111", 1 => "01101001", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            3059 => (0 => "01101001", 1 => "01101010", 2 => "01101011", 3 => "01101011", 4 => "11111111"),
            3060 => (0 => "11101100", 1 => "00101100", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            3061 => (0 => "00101100", 1 => "01001100", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            3062 => (0 => "01001100", 1 => "01111100", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            3063 => (0 => "01111100", 1 => "01100100", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            3064 => (0 => "01100100", 1 => "01101000", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            3065 => (0 => "01101000", 1 => "01101110", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            3066 => (0 => "01101110", 1 => "01101101", 2 => "01101100", 3 => "01101100", 4 => "11111111"),
            3067 => (0 => "11101101", 1 => "00101101", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            3068 => (0 => "00101101", 1 => "01001101", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            3069 => (0 => "01001101", 1 => "01111101", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            3070 => (0 => "01111101", 1 => "01100101", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            3071 => (0 => "01100101", 1 => "01101001", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            3072 => (0 => "01101001", 1 => "01101111", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            3073 => (0 => "01101111", 1 => "01101100", 2 => "01101101", 3 => "01101101", 4 => "11111111"),
            3074 => (0 => "11101110", 1 => "00101110", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            3075 => (0 => "00101110", 1 => "01001110", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            3076 => (0 => "01001110", 1 => "01111110", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            3077 => (0 => "01111110", 1 => "01100110", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            3078 => (0 => "01100110", 1 => "01101010", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            3079 => (0 => "01101010", 1 => "01101100", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            3080 => (0 => "01101100", 1 => "01101111", 2 => "01101110", 3 => "01101110", 4 => "11111111"),
            3081 => (0 => "11101111", 1 => "00101111", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            3082 => (0 => "00101111", 1 => "01001111", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            3083 => (0 => "01001111", 1 => "01111111", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            3084 => (0 => "01111111", 1 => "01100111", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            3085 => (0 => "01100111", 1 => "01101011", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            3086 => (0 => "01101011", 1 => "01101101", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            3087 => (0 => "01101101", 1 => "01101110", 2 => "01101111", 3 => "01101111", 4 => "11111111"),
            3088 => (0 => "11110000", 1 => "00110000", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            3089 => (0 => "00110000", 1 => "01010000", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            3090 => (0 => "01010000", 1 => "01100000", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            3091 => (0 => "01100000", 1 => "01111000", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            3092 => (0 => "01111000", 1 => "01110100", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            3093 => (0 => "01110100", 1 => "01110010", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            3094 => (0 => "01110010", 1 => "01110001", 2 => "01110000", 3 => "01110000", 4 => "11111111"),
            3095 => (0 => "11110001", 1 => "00110001", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            3096 => (0 => "00110001", 1 => "01010001", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            3097 => (0 => "01010001", 1 => "01100001", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            3098 => (0 => "01100001", 1 => "01111001", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            3099 => (0 => "01111001", 1 => "01110101", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            3100 => (0 => "01110101", 1 => "01110011", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            3101 => (0 => "01110011", 1 => "01110000", 2 => "01110001", 3 => "01110001", 4 => "11111111"),
            3102 => (0 => "11110010", 1 => "00110010", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            3103 => (0 => "00110010", 1 => "01010010", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            3104 => (0 => "01010010", 1 => "01100010", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            3105 => (0 => "01100010", 1 => "01111010", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            3106 => (0 => "01111010", 1 => "01110110", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            3107 => (0 => "01110110", 1 => "01110000", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            3108 => (0 => "01110000", 1 => "01110011", 2 => "01110010", 3 => "01110010", 4 => "11111111"),
            3109 => (0 => "11110011", 1 => "00110011", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            3110 => (0 => "00110011", 1 => "01010011", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            3111 => (0 => "01010011", 1 => "01100011", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            3112 => (0 => "01100011", 1 => "01111011", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            3113 => (0 => "01111011", 1 => "01110111", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            3114 => (0 => "01110111", 1 => "01110001", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            3115 => (0 => "01110001", 1 => "01110010", 2 => "01110011", 3 => "01110011", 4 => "11111111"),
            3116 => (0 => "11110100", 1 => "00110100", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            3117 => (0 => "00110100", 1 => "01010100", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            3118 => (0 => "01010100", 1 => "01100100", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            3119 => (0 => "01100100", 1 => "01111100", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            3120 => (0 => "01111100", 1 => "01110000", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            3121 => (0 => "01110000", 1 => "01110110", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            3122 => (0 => "01110110", 1 => "01110101", 2 => "01110100", 3 => "01110100", 4 => "11111111"),
            3123 => (0 => "11110101", 1 => "00110101", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            3124 => (0 => "00110101", 1 => "01010101", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            3125 => (0 => "01010101", 1 => "01100101", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            3126 => (0 => "01100101", 1 => "01111101", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            3127 => (0 => "01111101", 1 => "01110001", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            3128 => (0 => "01110001", 1 => "01110111", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            3129 => (0 => "01110111", 1 => "01110100", 2 => "01110101", 3 => "01110101", 4 => "11111111"),
            3130 => (0 => "11110110", 1 => "00110110", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            3131 => (0 => "00110110", 1 => "01010110", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            3132 => (0 => "01010110", 1 => "01100110", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            3133 => (0 => "01100110", 1 => "01111110", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            3134 => (0 => "01111110", 1 => "01110010", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            3135 => (0 => "01110010", 1 => "01110100", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            3136 => (0 => "01110100", 1 => "01110111", 2 => "01110110", 3 => "01110110", 4 => "11111111"),
            3137 => (0 => "11110111", 1 => "00110111", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            3138 => (0 => "00110111", 1 => "01010111", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            3139 => (0 => "01010111", 1 => "01100111", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            3140 => (0 => "01100111", 1 => "01111111", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            3141 => (0 => "01111111", 1 => "01110011", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            3142 => (0 => "01110011", 1 => "01110101", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            3143 => (0 => "01110101", 1 => "01110110", 2 => "01110111", 3 => "01110111", 4 => "11111111"),
            3144 => (0 => "11111000", 1 => "00111000", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            3145 => (0 => "00111000", 1 => "01011000", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            3146 => (0 => "01011000", 1 => "01101000", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            3147 => (0 => "01101000", 1 => "01110000", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            3148 => (0 => "01110000", 1 => "01111100", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            3149 => (0 => "01111100", 1 => "01111010", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            3150 => (0 => "01111010", 1 => "01111001", 2 => "01111000", 3 => "01111000", 4 => "11111111"),
            3151 => (0 => "11111001", 1 => "00111001", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            3152 => (0 => "00111001", 1 => "01011001", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            3153 => (0 => "01011001", 1 => "01101001", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            3154 => (0 => "01101001", 1 => "01110001", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            3155 => (0 => "01110001", 1 => "01111101", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            3156 => (0 => "01111101", 1 => "01111011", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            3157 => (0 => "01111011", 1 => "01111000", 2 => "01111001", 3 => "01111001", 4 => "11111111"),
            3158 => (0 => "11111010", 1 => "00111010", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            3159 => (0 => "00111010", 1 => "01011010", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            3160 => (0 => "01011010", 1 => "01101010", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            3161 => (0 => "01101010", 1 => "01110010", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            3162 => (0 => "01110010", 1 => "01111110", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            3163 => (0 => "01111110", 1 => "01111000", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            3164 => (0 => "01111000", 1 => "01111011", 2 => "01111010", 3 => "01111010", 4 => "11111111"),
            3165 => (0 => "11111011", 1 => "00111011", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            3166 => (0 => "00111011", 1 => "01011011", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            3167 => (0 => "01011011", 1 => "01101011", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            3168 => (0 => "01101011", 1 => "01110011", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            3169 => (0 => "01110011", 1 => "01111111", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            3170 => (0 => "01111111", 1 => "01111001", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            3171 => (0 => "01111001", 1 => "01111010", 2 => "01111011", 3 => "01111011", 4 => "11111111"),
            3172 => (0 => "11111100", 1 => "00111100", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            3173 => (0 => "00111100", 1 => "01011100", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            3174 => (0 => "01011100", 1 => "01101100", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            3175 => (0 => "01101100", 1 => "01110100", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            3176 => (0 => "01110100", 1 => "01111000", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            3177 => (0 => "01111000", 1 => "01111110", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            3178 => (0 => "01111110", 1 => "01111101", 2 => "01111100", 3 => "01111100", 4 => "11111111"),
            3179 => (0 => "11111101", 1 => "00111101", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            3180 => (0 => "00111101", 1 => "01011101", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            3181 => (0 => "01011101", 1 => "01101101", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            3182 => (0 => "01101101", 1 => "01110101", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            3183 => (0 => "01110101", 1 => "01111001", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            3184 => (0 => "01111001", 1 => "01111111", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            3185 => (0 => "01111111", 1 => "01111100", 2 => "01111101", 3 => "01111101", 4 => "11111111"),
            3186 => (0 => "11111110", 1 => "00111110", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            3187 => (0 => "00111110", 1 => "01011110", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            3188 => (0 => "01011110", 1 => "01101110", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            3189 => (0 => "01101110", 1 => "01110110", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            3190 => (0 => "01110110", 1 => "01111010", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            3191 => (0 => "01111010", 1 => "01111100", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            3192 => (0 => "01111100", 1 => "01111111", 2 => "01111110", 3 => "01111110", 4 => "11111111"),
            3193 => (0 => "11111111", 1 => "00111111", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            3194 => (0 => "00111111", 1 => "01011111", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            3195 => (0 => "01011111", 1 => "01101111", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            3196 => (0 => "01101111", 1 => "01110111", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            3197 => (0 => "01110111", 1 => "01111011", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            3198 => (0 => "01111011", 1 => "01111101", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            3199 => (0 => "01111101", 1 => "01111110", 2 => "01111111", 3 => "01111111", 4 => "11111111"),
            3200 => (0 => "00000000", 1 => "11000000", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            3201 => (0 => "11000000", 1 => "10100000", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            3202 => (0 => "10100000", 1 => "10010000", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            3203 => (0 => "10010000", 1 => "10001000", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            3204 => (0 => "10001000", 1 => "10000100", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            3205 => (0 => "10000100", 1 => "10000010", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            3206 => (0 => "10000010", 1 => "10000001", 2 => "10000000", 3 => "10000000", 4 => "11111111"),
            3207 => (0 => "00000001", 1 => "11000001", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            3208 => (0 => "11000001", 1 => "10100001", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            3209 => (0 => "10100001", 1 => "10010001", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            3210 => (0 => "10010001", 1 => "10001001", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            3211 => (0 => "10001001", 1 => "10000101", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            3212 => (0 => "10000101", 1 => "10000011", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            3213 => (0 => "10000011", 1 => "10000000", 2 => "10000001", 3 => "10000001", 4 => "11111111"),
            3214 => (0 => "00000010", 1 => "11000010", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            3215 => (0 => "11000010", 1 => "10100010", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            3216 => (0 => "10100010", 1 => "10010010", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            3217 => (0 => "10010010", 1 => "10001010", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            3218 => (0 => "10001010", 1 => "10000110", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            3219 => (0 => "10000110", 1 => "10000000", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            3220 => (0 => "10000000", 1 => "10000011", 2 => "10000010", 3 => "10000010", 4 => "11111111"),
            3221 => (0 => "00000011", 1 => "11000011", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            3222 => (0 => "11000011", 1 => "10100011", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            3223 => (0 => "10100011", 1 => "10010011", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            3224 => (0 => "10010011", 1 => "10001011", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            3225 => (0 => "10001011", 1 => "10000111", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            3226 => (0 => "10000111", 1 => "10000001", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            3227 => (0 => "10000001", 1 => "10000010", 2 => "10000011", 3 => "10000011", 4 => "11111111"),
            3228 => (0 => "00000100", 1 => "11000100", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            3229 => (0 => "11000100", 1 => "10100100", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            3230 => (0 => "10100100", 1 => "10010100", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            3231 => (0 => "10010100", 1 => "10001100", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            3232 => (0 => "10001100", 1 => "10000000", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            3233 => (0 => "10000000", 1 => "10000110", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            3234 => (0 => "10000110", 1 => "10000101", 2 => "10000100", 3 => "10000100", 4 => "11111111"),
            3235 => (0 => "00000101", 1 => "11000101", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            3236 => (0 => "11000101", 1 => "10100101", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            3237 => (0 => "10100101", 1 => "10010101", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            3238 => (0 => "10010101", 1 => "10001101", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            3239 => (0 => "10001101", 1 => "10000001", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            3240 => (0 => "10000001", 1 => "10000111", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            3241 => (0 => "10000111", 1 => "10000100", 2 => "10000101", 3 => "10000101", 4 => "11111111"),
            3242 => (0 => "00000110", 1 => "11000110", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            3243 => (0 => "11000110", 1 => "10100110", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            3244 => (0 => "10100110", 1 => "10010110", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            3245 => (0 => "10010110", 1 => "10001110", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            3246 => (0 => "10001110", 1 => "10000010", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            3247 => (0 => "10000010", 1 => "10000100", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            3248 => (0 => "10000100", 1 => "10000111", 2 => "10000110", 3 => "10000110", 4 => "11111111"),
            3249 => (0 => "00000111", 1 => "11000111", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            3250 => (0 => "11000111", 1 => "10100111", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            3251 => (0 => "10100111", 1 => "10010111", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            3252 => (0 => "10010111", 1 => "10001111", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            3253 => (0 => "10001111", 1 => "10000011", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            3254 => (0 => "10000011", 1 => "10000101", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            3255 => (0 => "10000101", 1 => "10000110", 2 => "10000111", 3 => "10000111", 4 => "11111111"),
            3256 => (0 => "00001000", 1 => "11001000", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            3257 => (0 => "11001000", 1 => "10101000", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            3258 => (0 => "10101000", 1 => "10011000", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            3259 => (0 => "10011000", 1 => "10000000", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            3260 => (0 => "10000000", 1 => "10001100", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            3261 => (0 => "10001100", 1 => "10001010", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            3262 => (0 => "10001010", 1 => "10001001", 2 => "10001000", 3 => "10001000", 4 => "11111111"),
            3263 => (0 => "00001001", 1 => "11001001", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            3264 => (0 => "11001001", 1 => "10101001", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            3265 => (0 => "10101001", 1 => "10011001", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            3266 => (0 => "10011001", 1 => "10000001", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            3267 => (0 => "10000001", 1 => "10001101", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            3268 => (0 => "10001101", 1 => "10001011", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            3269 => (0 => "10001011", 1 => "10001000", 2 => "10001001", 3 => "10001001", 4 => "11111111"),
            3270 => (0 => "00001010", 1 => "11001010", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            3271 => (0 => "11001010", 1 => "10101010", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            3272 => (0 => "10101010", 1 => "10011010", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            3273 => (0 => "10011010", 1 => "10000010", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            3274 => (0 => "10000010", 1 => "10001110", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            3275 => (0 => "10001110", 1 => "10001000", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            3276 => (0 => "10001000", 1 => "10001011", 2 => "10001010", 3 => "10001010", 4 => "11111111"),
            3277 => (0 => "00001011", 1 => "11001011", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            3278 => (0 => "11001011", 1 => "10101011", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            3279 => (0 => "10101011", 1 => "10011011", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            3280 => (0 => "10011011", 1 => "10000011", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            3281 => (0 => "10000011", 1 => "10001111", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            3282 => (0 => "10001111", 1 => "10001001", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            3283 => (0 => "10001001", 1 => "10001010", 2 => "10001011", 3 => "10001011", 4 => "11111111"),
            3284 => (0 => "00001100", 1 => "11001100", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            3285 => (0 => "11001100", 1 => "10101100", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            3286 => (0 => "10101100", 1 => "10011100", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            3287 => (0 => "10011100", 1 => "10000100", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            3288 => (0 => "10000100", 1 => "10001000", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            3289 => (0 => "10001000", 1 => "10001110", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            3290 => (0 => "10001110", 1 => "10001101", 2 => "10001100", 3 => "10001100", 4 => "11111111"),
            3291 => (0 => "00001101", 1 => "11001101", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            3292 => (0 => "11001101", 1 => "10101101", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            3293 => (0 => "10101101", 1 => "10011101", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            3294 => (0 => "10011101", 1 => "10000101", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            3295 => (0 => "10000101", 1 => "10001001", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            3296 => (0 => "10001001", 1 => "10001111", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            3297 => (0 => "10001111", 1 => "10001100", 2 => "10001101", 3 => "10001101", 4 => "11111111"),
            3298 => (0 => "00001110", 1 => "11001110", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            3299 => (0 => "11001110", 1 => "10101110", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            3300 => (0 => "10101110", 1 => "10011110", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            3301 => (0 => "10011110", 1 => "10000110", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            3302 => (0 => "10000110", 1 => "10001010", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            3303 => (0 => "10001010", 1 => "10001100", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            3304 => (0 => "10001100", 1 => "10001111", 2 => "10001110", 3 => "10001110", 4 => "11111111"),
            3305 => (0 => "00001111", 1 => "11001111", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            3306 => (0 => "11001111", 1 => "10101111", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            3307 => (0 => "10101111", 1 => "10011111", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            3308 => (0 => "10011111", 1 => "10000111", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            3309 => (0 => "10000111", 1 => "10001011", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            3310 => (0 => "10001011", 1 => "10001101", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            3311 => (0 => "10001101", 1 => "10001110", 2 => "10001111", 3 => "10001111", 4 => "11111111"),
            3312 => (0 => "00010000", 1 => "11010000", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            3313 => (0 => "11010000", 1 => "10110000", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            3314 => (0 => "10110000", 1 => "10000000", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            3315 => (0 => "10000000", 1 => "10011000", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            3316 => (0 => "10011000", 1 => "10010100", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            3317 => (0 => "10010100", 1 => "10010010", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            3318 => (0 => "10010010", 1 => "10010001", 2 => "10010000", 3 => "10010000", 4 => "11111111"),
            3319 => (0 => "00010001", 1 => "11010001", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            3320 => (0 => "11010001", 1 => "10110001", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            3321 => (0 => "10110001", 1 => "10000001", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            3322 => (0 => "10000001", 1 => "10011001", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            3323 => (0 => "10011001", 1 => "10010101", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            3324 => (0 => "10010101", 1 => "10010011", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            3325 => (0 => "10010011", 1 => "10010000", 2 => "10010001", 3 => "10010001", 4 => "11111111"),
            3326 => (0 => "00010010", 1 => "11010010", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            3327 => (0 => "11010010", 1 => "10110010", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            3328 => (0 => "10110010", 1 => "10000010", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            3329 => (0 => "10000010", 1 => "10011010", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            3330 => (0 => "10011010", 1 => "10010110", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            3331 => (0 => "10010110", 1 => "10010000", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            3332 => (0 => "10010000", 1 => "10010011", 2 => "10010010", 3 => "10010010", 4 => "11111111"),
            3333 => (0 => "00010011", 1 => "11010011", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            3334 => (0 => "11010011", 1 => "10110011", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            3335 => (0 => "10110011", 1 => "10000011", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            3336 => (0 => "10000011", 1 => "10011011", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            3337 => (0 => "10011011", 1 => "10010111", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            3338 => (0 => "10010111", 1 => "10010001", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            3339 => (0 => "10010001", 1 => "10010010", 2 => "10010011", 3 => "10010011", 4 => "11111111"),
            3340 => (0 => "00010100", 1 => "11010100", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            3341 => (0 => "11010100", 1 => "10110100", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            3342 => (0 => "10110100", 1 => "10000100", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            3343 => (0 => "10000100", 1 => "10011100", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            3344 => (0 => "10011100", 1 => "10010000", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            3345 => (0 => "10010000", 1 => "10010110", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            3346 => (0 => "10010110", 1 => "10010101", 2 => "10010100", 3 => "10010100", 4 => "11111111"),
            3347 => (0 => "00010101", 1 => "11010101", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            3348 => (0 => "11010101", 1 => "10110101", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            3349 => (0 => "10110101", 1 => "10000101", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            3350 => (0 => "10000101", 1 => "10011101", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            3351 => (0 => "10011101", 1 => "10010001", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            3352 => (0 => "10010001", 1 => "10010111", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            3353 => (0 => "10010111", 1 => "10010100", 2 => "10010101", 3 => "10010101", 4 => "11111111"),
            3354 => (0 => "00010110", 1 => "11010110", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            3355 => (0 => "11010110", 1 => "10110110", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            3356 => (0 => "10110110", 1 => "10000110", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            3357 => (0 => "10000110", 1 => "10011110", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            3358 => (0 => "10011110", 1 => "10010010", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            3359 => (0 => "10010010", 1 => "10010100", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            3360 => (0 => "10010100", 1 => "10010111", 2 => "10010110", 3 => "10010110", 4 => "11111111"),
            3361 => (0 => "00010111", 1 => "11010111", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            3362 => (0 => "11010111", 1 => "10110111", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            3363 => (0 => "10110111", 1 => "10000111", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            3364 => (0 => "10000111", 1 => "10011111", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            3365 => (0 => "10011111", 1 => "10010011", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            3366 => (0 => "10010011", 1 => "10010101", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            3367 => (0 => "10010101", 1 => "10010110", 2 => "10010111", 3 => "10010111", 4 => "11111111"),
            3368 => (0 => "00011000", 1 => "11011000", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            3369 => (0 => "11011000", 1 => "10111000", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            3370 => (0 => "10111000", 1 => "10001000", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            3371 => (0 => "10001000", 1 => "10010000", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            3372 => (0 => "10010000", 1 => "10011100", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            3373 => (0 => "10011100", 1 => "10011010", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            3374 => (0 => "10011010", 1 => "10011001", 2 => "10011000", 3 => "10011000", 4 => "11111111"),
            3375 => (0 => "00011001", 1 => "11011001", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            3376 => (0 => "11011001", 1 => "10111001", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            3377 => (0 => "10111001", 1 => "10001001", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            3378 => (0 => "10001001", 1 => "10010001", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            3379 => (0 => "10010001", 1 => "10011101", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            3380 => (0 => "10011101", 1 => "10011011", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            3381 => (0 => "10011011", 1 => "10011000", 2 => "10011001", 3 => "10011001", 4 => "11111111"),
            3382 => (0 => "00011010", 1 => "11011010", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            3383 => (0 => "11011010", 1 => "10111010", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            3384 => (0 => "10111010", 1 => "10001010", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            3385 => (0 => "10001010", 1 => "10010010", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            3386 => (0 => "10010010", 1 => "10011110", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            3387 => (0 => "10011110", 1 => "10011000", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            3388 => (0 => "10011000", 1 => "10011011", 2 => "10011010", 3 => "10011010", 4 => "11111111"),
            3389 => (0 => "00011011", 1 => "11011011", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            3390 => (0 => "11011011", 1 => "10111011", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            3391 => (0 => "10111011", 1 => "10001011", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            3392 => (0 => "10001011", 1 => "10010011", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            3393 => (0 => "10010011", 1 => "10011111", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            3394 => (0 => "10011111", 1 => "10011001", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            3395 => (0 => "10011001", 1 => "10011010", 2 => "10011011", 3 => "10011011", 4 => "11111111"),
            3396 => (0 => "00011100", 1 => "11011100", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            3397 => (0 => "11011100", 1 => "10111100", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            3398 => (0 => "10111100", 1 => "10001100", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            3399 => (0 => "10001100", 1 => "10010100", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            3400 => (0 => "10010100", 1 => "10011000", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            3401 => (0 => "10011000", 1 => "10011110", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            3402 => (0 => "10011110", 1 => "10011101", 2 => "10011100", 3 => "10011100", 4 => "11111111"),
            3403 => (0 => "00011101", 1 => "11011101", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            3404 => (0 => "11011101", 1 => "10111101", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            3405 => (0 => "10111101", 1 => "10001101", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            3406 => (0 => "10001101", 1 => "10010101", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            3407 => (0 => "10010101", 1 => "10011001", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            3408 => (0 => "10011001", 1 => "10011111", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            3409 => (0 => "10011111", 1 => "10011100", 2 => "10011101", 3 => "10011101", 4 => "11111111"),
            3410 => (0 => "00011110", 1 => "11011110", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            3411 => (0 => "11011110", 1 => "10111110", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            3412 => (0 => "10111110", 1 => "10001110", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            3413 => (0 => "10001110", 1 => "10010110", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            3414 => (0 => "10010110", 1 => "10011010", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            3415 => (0 => "10011010", 1 => "10011100", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            3416 => (0 => "10011100", 1 => "10011111", 2 => "10011110", 3 => "10011110", 4 => "11111111"),
            3417 => (0 => "00011111", 1 => "11011111", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            3418 => (0 => "11011111", 1 => "10111111", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            3419 => (0 => "10111111", 1 => "10001111", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            3420 => (0 => "10001111", 1 => "10010111", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            3421 => (0 => "10010111", 1 => "10011011", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            3422 => (0 => "10011011", 1 => "10011101", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            3423 => (0 => "10011101", 1 => "10011110", 2 => "10011111", 3 => "10011111", 4 => "11111111"),
            3424 => (0 => "00100000", 1 => "11100000", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            3425 => (0 => "11100000", 1 => "10000000", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            3426 => (0 => "10000000", 1 => "10110000", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            3427 => (0 => "10110000", 1 => "10101000", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            3428 => (0 => "10101000", 1 => "10100100", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            3429 => (0 => "10100100", 1 => "10100010", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            3430 => (0 => "10100010", 1 => "10100001", 2 => "10100000", 3 => "10100000", 4 => "11111111"),
            3431 => (0 => "00100001", 1 => "11100001", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            3432 => (0 => "11100001", 1 => "10000001", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            3433 => (0 => "10000001", 1 => "10110001", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            3434 => (0 => "10110001", 1 => "10101001", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            3435 => (0 => "10101001", 1 => "10100101", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            3436 => (0 => "10100101", 1 => "10100011", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            3437 => (0 => "10100011", 1 => "10100000", 2 => "10100001", 3 => "10100001", 4 => "11111111"),
            3438 => (0 => "00100010", 1 => "11100010", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            3439 => (0 => "11100010", 1 => "10000010", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            3440 => (0 => "10000010", 1 => "10110010", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            3441 => (0 => "10110010", 1 => "10101010", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            3442 => (0 => "10101010", 1 => "10100110", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            3443 => (0 => "10100110", 1 => "10100000", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            3444 => (0 => "10100000", 1 => "10100011", 2 => "10100010", 3 => "10100010", 4 => "11111111"),
            3445 => (0 => "00100011", 1 => "11100011", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            3446 => (0 => "11100011", 1 => "10000011", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            3447 => (0 => "10000011", 1 => "10110011", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            3448 => (0 => "10110011", 1 => "10101011", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            3449 => (0 => "10101011", 1 => "10100111", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            3450 => (0 => "10100111", 1 => "10100001", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            3451 => (0 => "10100001", 1 => "10100010", 2 => "10100011", 3 => "10100011", 4 => "11111111"),
            3452 => (0 => "00100100", 1 => "11100100", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            3453 => (0 => "11100100", 1 => "10000100", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            3454 => (0 => "10000100", 1 => "10110100", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            3455 => (0 => "10110100", 1 => "10101100", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            3456 => (0 => "10101100", 1 => "10100000", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            3457 => (0 => "10100000", 1 => "10100110", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            3458 => (0 => "10100110", 1 => "10100101", 2 => "10100100", 3 => "10100100", 4 => "11111111"),
            3459 => (0 => "00100101", 1 => "11100101", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            3460 => (0 => "11100101", 1 => "10000101", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            3461 => (0 => "10000101", 1 => "10110101", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            3462 => (0 => "10110101", 1 => "10101101", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            3463 => (0 => "10101101", 1 => "10100001", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            3464 => (0 => "10100001", 1 => "10100111", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            3465 => (0 => "10100111", 1 => "10100100", 2 => "10100101", 3 => "10100101", 4 => "11111111"),
            3466 => (0 => "00100110", 1 => "11100110", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            3467 => (0 => "11100110", 1 => "10000110", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            3468 => (0 => "10000110", 1 => "10110110", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            3469 => (0 => "10110110", 1 => "10101110", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            3470 => (0 => "10101110", 1 => "10100010", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            3471 => (0 => "10100010", 1 => "10100100", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            3472 => (0 => "10100100", 1 => "10100111", 2 => "10100110", 3 => "10100110", 4 => "11111111"),
            3473 => (0 => "00100111", 1 => "11100111", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            3474 => (0 => "11100111", 1 => "10000111", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            3475 => (0 => "10000111", 1 => "10110111", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            3476 => (0 => "10110111", 1 => "10101111", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            3477 => (0 => "10101111", 1 => "10100011", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            3478 => (0 => "10100011", 1 => "10100101", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            3479 => (0 => "10100101", 1 => "10100110", 2 => "10100111", 3 => "10100111", 4 => "11111111"),
            3480 => (0 => "00101000", 1 => "11101000", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            3481 => (0 => "11101000", 1 => "10001000", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            3482 => (0 => "10001000", 1 => "10111000", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            3483 => (0 => "10111000", 1 => "10100000", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            3484 => (0 => "10100000", 1 => "10101100", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            3485 => (0 => "10101100", 1 => "10101010", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            3486 => (0 => "10101010", 1 => "10101001", 2 => "10101000", 3 => "10101000", 4 => "11111111"),
            3487 => (0 => "00101001", 1 => "11101001", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            3488 => (0 => "11101001", 1 => "10001001", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            3489 => (0 => "10001001", 1 => "10111001", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            3490 => (0 => "10111001", 1 => "10100001", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            3491 => (0 => "10100001", 1 => "10101101", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            3492 => (0 => "10101101", 1 => "10101011", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            3493 => (0 => "10101011", 1 => "10101000", 2 => "10101001", 3 => "10101001", 4 => "11111111"),
            3494 => (0 => "00101010", 1 => "11101010", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            3495 => (0 => "11101010", 1 => "10001010", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            3496 => (0 => "10001010", 1 => "10111010", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            3497 => (0 => "10111010", 1 => "10100010", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            3498 => (0 => "10100010", 1 => "10101110", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            3499 => (0 => "10101110", 1 => "10101000", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            3500 => (0 => "10101000", 1 => "10101011", 2 => "10101010", 3 => "10101010", 4 => "11111111"),
            3501 => (0 => "00101011", 1 => "11101011", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            3502 => (0 => "11101011", 1 => "10001011", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            3503 => (0 => "10001011", 1 => "10111011", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            3504 => (0 => "10111011", 1 => "10100011", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            3505 => (0 => "10100011", 1 => "10101111", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            3506 => (0 => "10101111", 1 => "10101001", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            3507 => (0 => "10101001", 1 => "10101010", 2 => "10101011", 3 => "10101011", 4 => "11111111"),
            3508 => (0 => "00101100", 1 => "11101100", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            3509 => (0 => "11101100", 1 => "10001100", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            3510 => (0 => "10001100", 1 => "10111100", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            3511 => (0 => "10111100", 1 => "10100100", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            3512 => (0 => "10100100", 1 => "10101000", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            3513 => (0 => "10101000", 1 => "10101110", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            3514 => (0 => "10101110", 1 => "10101101", 2 => "10101100", 3 => "10101100", 4 => "11111111"),
            3515 => (0 => "00101101", 1 => "11101101", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            3516 => (0 => "11101101", 1 => "10001101", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            3517 => (0 => "10001101", 1 => "10111101", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            3518 => (0 => "10111101", 1 => "10100101", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            3519 => (0 => "10100101", 1 => "10101001", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            3520 => (0 => "10101001", 1 => "10101111", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            3521 => (0 => "10101111", 1 => "10101100", 2 => "10101101", 3 => "10101101", 4 => "11111111"),
            3522 => (0 => "00101110", 1 => "11101110", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            3523 => (0 => "11101110", 1 => "10001110", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            3524 => (0 => "10001110", 1 => "10111110", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            3525 => (0 => "10111110", 1 => "10100110", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            3526 => (0 => "10100110", 1 => "10101010", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            3527 => (0 => "10101010", 1 => "10101100", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            3528 => (0 => "10101100", 1 => "10101111", 2 => "10101110", 3 => "10101110", 4 => "11111111"),
            3529 => (0 => "00101111", 1 => "11101111", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            3530 => (0 => "11101111", 1 => "10001111", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            3531 => (0 => "10001111", 1 => "10111111", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            3532 => (0 => "10111111", 1 => "10100111", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            3533 => (0 => "10100111", 1 => "10101011", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            3534 => (0 => "10101011", 1 => "10101101", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            3535 => (0 => "10101101", 1 => "10101110", 2 => "10101111", 3 => "10101111", 4 => "11111111"),
            3536 => (0 => "00110000", 1 => "11110000", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            3537 => (0 => "11110000", 1 => "10010000", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            3538 => (0 => "10010000", 1 => "10100000", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            3539 => (0 => "10100000", 1 => "10111000", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            3540 => (0 => "10111000", 1 => "10110100", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            3541 => (0 => "10110100", 1 => "10110010", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            3542 => (0 => "10110010", 1 => "10110001", 2 => "10110000", 3 => "10110000", 4 => "11111111"),
            3543 => (0 => "00110001", 1 => "11110001", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            3544 => (0 => "11110001", 1 => "10010001", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            3545 => (0 => "10010001", 1 => "10100001", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            3546 => (0 => "10100001", 1 => "10111001", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            3547 => (0 => "10111001", 1 => "10110101", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            3548 => (0 => "10110101", 1 => "10110011", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            3549 => (0 => "10110011", 1 => "10110000", 2 => "10110001", 3 => "10110001", 4 => "11111111"),
            3550 => (0 => "00110010", 1 => "11110010", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            3551 => (0 => "11110010", 1 => "10010010", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            3552 => (0 => "10010010", 1 => "10100010", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            3553 => (0 => "10100010", 1 => "10111010", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            3554 => (0 => "10111010", 1 => "10110110", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            3555 => (0 => "10110110", 1 => "10110000", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            3556 => (0 => "10110000", 1 => "10110011", 2 => "10110010", 3 => "10110010", 4 => "11111111"),
            3557 => (0 => "00110011", 1 => "11110011", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            3558 => (0 => "11110011", 1 => "10010011", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            3559 => (0 => "10010011", 1 => "10100011", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            3560 => (0 => "10100011", 1 => "10111011", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            3561 => (0 => "10111011", 1 => "10110111", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            3562 => (0 => "10110111", 1 => "10110001", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            3563 => (0 => "10110001", 1 => "10110010", 2 => "10110011", 3 => "10110011", 4 => "11111111"),
            3564 => (0 => "00110100", 1 => "11110100", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            3565 => (0 => "11110100", 1 => "10010100", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            3566 => (0 => "10010100", 1 => "10100100", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            3567 => (0 => "10100100", 1 => "10111100", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            3568 => (0 => "10111100", 1 => "10110000", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            3569 => (0 => "10110000", 1 => "10110110", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            3570 => (0 => "10110110", 1 => "10110101", 2 => "10110100", 3 => "10110100", 4 => "11111111"),
            3571 => (0 => "00110101", 1 => "11110101", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            3572 => (0 => "11110101", 1 => "10010101", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            3573 => (0 => "10010101", 1 => "10100101", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            3574 => (0 => "10100101", 1 => "10111101", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            3575 => (0 => "10111101", 1 => "10110001", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            3576 => (0 => "10110001", 1 => "10110111", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            3577 => (0 => "10110111", 1 => "10110100", 2 => "10110101", 3 => "10110101", 4 => "11111111"),
            3578 => (0 => "00110110", 1 => "11110110", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            3579 => (0 => "11110110", 1 => "10010110", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            3580 => (0 => "10010110", 1 => "10100110", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            3581 => (0 => "10100110", 1 => "10111110", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            3582 => (0 => "10111110", 1 => "10110010", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            3583 => (0 => "10110010", 1 => "10110100", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            3584 => (0 => "10110100", 1 => "10110111", 2 => "10110110", 3 => "10110110", 4 => "11111111"),
            3585 => (0 => "00110111", 1 => "11110111", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            3586 => (0 => "11110111", 1 => "10010111", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            3587 => (0 => "10010111", 1 => "10100111", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            3588 => (0 => "10100111", 1 => "10111111", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            3589 => (0 => "10111111", 1 => "10110011", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            3590 => (0 => "10110011", 1 => "10110101", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            3591 => (0 => "10110101", 1 => "10110110", 2 => "10110111", 3 => "10110111", 4 => "11111111"),
            3592 => (0 => "00111000", 1 => "11111000", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            3593 => (0 => "11111000", 1 => "10011000", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            3594 => (0 => "10011000", 1 => "10101000", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            3595 => (0 => "10101000", 1 => "10110000", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            3596 => (0 => "10110000", 1 => "10111100", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            3597 => (0 => "10111100", 1 => "10111010", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            3598 => (0 => "10111010", 1 => "10111001", 2 => "10111000", 3 => "10111000", 4 => "11111111"),
            3599 => (0 => "00111001", 1 => "11111001", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            3600 => (0 => "11111001", 1 => "10011001", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            3601 => (0 => "10011001", 1 => "10101001", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            3602 => (0 => "10101001", 1 => "10110001", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            3603 => (0 => "10110001", 1 => "10111101", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            3604 => (0 => "10111101", 1 => "10111011", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            3605 => (0 => "10111011", 1 => "10111000", 2 => "10111001", 3 => "10111001", 4 => "11111111"),
            3606 => (0 => "00111010", 1 => "11111010", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            3607 => (0 => "11111010", 1 => "10011010", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            3608 => (0 => "10011010", 1 => "10101010", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            3609 => (0 => "10101010", 1 => "10110010", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            3610 => (0 => "10110010", 1 => "10111110", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            3611 => (0 => "10111110", 1 => "10111000", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            3612 => (0 => "10111000", 1 => "10111011", 2 => "10111010", 3 => "10111010", 4 => "11111111"),
            3613 => (0 => "00111011", 1 => "11111011", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            3614 => (0 => "11111011", 1 => "10011011", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            3615 => (0 => "10011011", 1 => "10101011", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            3616 => (0 => "10101011", 1 => "10110011", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            3617 => (0 => "10110011", 1 => "10111111", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            3618 => (0 => "10111111", 1 => "10111001", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            3619 => (0 => "10111001", 1 => "10111010", 2 => "10111011", 3 => "10111011", 4 => "11111111"),
            3620 => (0 => "00111100", 1 => "11111100", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            3621 => (0 => "11111100", 1 => "10011100", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            3622 => (0 => "10011100", 1 => "10101100", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            3623 => (0 => "10101100", 1 => "10110100", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            3624 => (0 => "10110100", 1 => "10111000", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            3625 => (0 => "10111000", 1 => "10111110", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            3626 => (0 => "10111110", 1 => "10111101", 2 => "10111100", 3 => "10111100", 4 => "11111111"),
            3627 => (0 => "00111101", 1 => "11111101", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            3628 => (0 => "11111101", 1 => "10011101", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            3629 => (0 => "10011101", 1 => "10101101", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            3630 => (0 => "10101101", 1 => "10110101", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            3631 => (0 => "10110101", 1 => "10111001", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            3632 => (0 => "10111001", 1 => "10111111", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            3633 => (0 => "10111111", 1 => "10111100", 2 => "10111101", 3 => "10111101", 4 => "11111111"),
            3634 => (0 => "00111110", 1 => "11111110", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            3635 => (0 => "11111110", 1 => "10011110", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            3636 => (0 => "10011110", 1 => "10101110", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            3637 => (0 => "10101110", 1 => "10110110", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            3638 => (0 => "10110110", 1 => "10111010", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            3639 => (0 => "10111010", 1 => "10111100", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            3640 => (0 => "10111100", 1 => "10111111", 2 => "10111110", 3 => "10111110", 4 => "11111111"),
            3641 => (0 => "00111111", 1 => "11111111", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            3642 => (0 => "11111111", 1 => "10011111", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            3643 => (0 => "10011111", 1 => "10101111", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            3644 => (0 => "10101111", 1 => "10110111", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            3645 => (0 => "10110111", 1 => "10111011", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            3646 => (0 => "10111011", 1 => "10111101", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            3647 => (0 => "10111101", 1 => "10111110", 2 => "10111111", 3 => "10111111", 4 => "11111111"),
            3648 => (0 => "01000000", 1 => "10000000", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            3649 => (0 => "10000000", 1 => "11100000", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            3650 => (0 => "11100000", 1 => "11010000", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            3651 => (0 => "11010000", 1 => "11001000", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            3652 => (0 => "11001000", 1 => "11000100", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            3653 => (0 => "11000100", 1 => "11000010", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            3654 => (0 => "11000010", 1 => "11000001", 2 => "11000000", 3 => "11000000", 4 => "11111111"),
            3655 => (0 => "01000001", 1 => "10000001", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            3656 => (0 => "10000001", 1 => "11100001", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            3657 => (0 => "11100001", 1 => "11010001", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            3658 => (0 => "11010001", 1 => "11001001", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            3659 => (0 => "11001001", 1 => "11000101", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            3660 => (0 => "11000101", 1 => "11000011", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            3661 => (0 => "11000011", 1 => "11000000", 2 => "11000001", 3 => "11000001", 4 => "11111111"),
            3662 => (0 => "01000010", 1 => "10000010", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            3663 => (0 => "10000010", 1 => "11100010", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            3664 => (0 => "11100010", 1 => "11010010", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            3665 => (0 => "11010010", 1 => "11001010", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            3666 => (0 => "11001010", 1 => "11000110", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            3667 => (0 => "11000110", 1 => "11000000", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            3668 => (0 => "11000000", 1 => "11000011", 2 => "11000010", 3 => "11000010", 4 => "11111111"),
            3669 => (0 => "01000011", 1 => "10000011", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            3670 => (0 => "10000011", 1 => "11100011", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            3671 => (0 => "11100011", 1 => "11010011", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            3672 => (0 => "11010011", 1 => "11001011", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            3673 => (0 => "11001011", 1 => "11000111", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            3674 => (0 => "11000111", 1 => "11000001", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            3675 => (0 => "11000001", 1 => "11000010", 2 => "11000011", 3 => "11000011", 4 => "11111111"),
            3676 => (0 => "01000100", 1 => "10000100", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            3677 => (0 => "10000100", 1 => "11100100", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            3678 => (0 => "11100100", 1 => "11010100", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            3679 => (0 => "11010100", 1 => "11001100", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            3680 => (0 => "11001100", 1 => "11000000", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            3681 => (0 => "11000000", 1 => "11000110", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            3682 => (0 => "11000110", 1 => "11000101", 2 => "11000100", 3 => "11000100", 4 => "11111111"),
            3683 => (0 => "01000101", 1 => "10000101", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            3684 => (0 => "10000101", 1 => "11100101", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            3685 => (0 => "11100101", 1 => "11010101", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            3686 => (0 => "11010101", 1 => "11001101", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            3687 => (0 => "11001101", 1 => "11000001", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            3688 => (0 => "11000001", 1 => "11000111", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            3689 => (0 => "11000111", 1 => "11000100", 2 => "11000101", 3 => "11000101", 4 => "11111111"),
            3690 => (0 => "01000110", 1 => "10000110", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            3691 => (0 => "10000110", 1 => "11100110", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            3692 => (0 => "11100110", 1 => "11010110", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            3693 => (0 => "11010110", 1 => "11001110", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            3694 => (0 => "11001110", 1 => "11000010", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            3695 => (0 => "11000010", 1 => "11000100", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            3696 => (0 => "11000100", 1 => "11000111", 2 => "11000110", 3 => "11000110", 4 => "11111111"),
            3697 => (0 => "01000111", 1 => "10000111", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            3698 => (0 => "10000111", 1 => "11100111", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            3699 => (0 => "11100111", 1 => "11010111", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            3700 => (0 => "11010111", 1 => "11001111", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            3701 => (0 => "11001111", 1 => "11000011", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            3702 => (0 => "11000011", 1 => "11000101", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            3703 => (0 => "11000101", 1 => "11000110", 2 => "11000111", 3 => "11000111", 4 => "11111111"),
            3704 => (0 => "01001000", 1 => "10001000", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            3705 => (0 => "10001000", 1 => "11101000", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            3706 => (0 => "11101000", 1 => "11011000", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            3707 => (0 => "11011000", 1 => "11000000", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            3708 => (0 => "11000000", 1 => "11001100", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            3709 => (0 => "11001100", 1 => "11001010", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            3710 => (0 => "11001010", 1 => "11001001", 2 => "11001000", 3 => "11001000", 4 => "11111111"),
            3711 => (0 => "01001001", 1 => "10001001", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            3712 => (0 => "10001001", 1 => "11101001", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            3713 => (0 => "11101001", 1 => "11011001", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            3714 => (0 => "11011001", 1 => "11000001", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            3715 => (0 => "11000001", 1 => "11001101", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            3716 => (0 => "11001101", 1 => "11001011", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            3717 => (0 => "11001011", 1 => "11001000", 2 => "11001001", 3 => "11001001", 4 => "11111111"),
            3718 => (0 => "01001010", 1 => "10001010", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            3719 => (0 => "10001010", 1 => "11101010", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            3720 => (0 => "11101010", 1 => "11011010", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            3721 => (0 => "11011010", 1 => "11000010", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            3722 => (0 => "11000010", 1 => "11001110", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            3723 => (0 => "11001110", 1 => "11001000", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            3724 => (0 => "11001000", 1 => "11001011", 2 => "11001010", 3 => "11001010", 4 => "11111111"),
            3725 => (0 => "01001011", 1 => "10001011", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            3726 => (0 => "10001011", 1 => "11101011", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            3727 => (0 => "11101011", 1 => "11011011", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            3728 => (0 => "11011011", 1 => "11000011", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            3729 => (0 => "11000011", 1 => "11001111", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            3730 => (0 => "11001111", 1 => "11001001", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            3731 => (0 => "11001001", 1 => "11001010", 2 => "11001011", 3 => "11001011", 4 => "11111111"),
            3732 => (0 => "01001100", 1 => "10001100", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            3733 => (0 => "10001100", 1 => "11101100", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            3734 => (0 => "11101100", 1 => "11011100", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            3735 => (0 => "11011100", 1 => "11000100", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            3736 => (0 => "11000100", 1 => "11001000", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            3737 => (0 => "11001000", 1 => "11001110", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            3738 => (0 => "11001110", 1 => "11001101", 2 => "11001100", 3 => "11001100", 4 => "11111111"),
            3739 => (0 => "01001101", 1 => "10001101", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            3740 => (0 => "10001101", 1 => "11101101", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            3741 => (0 => "11101101", 1 => "11011101", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            3742 => (0 => "11011101", 1 => "11000101", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            3743 => (0 => "11000101", 1 => "11001001", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            3744 => (0 => "11001001", 1 => "11001111", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            3745 => (0 => "11001111", 1 => "11001100", 2 => "11001101", 3 => "11001101", 4 => "11111111"),
            3746 => (0 => "01001110", 1 => "10001110", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            3747 => (0 => "10001110", 1 => "11101110", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            3748 => (0 => "11101110", 1 => "11011110", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            3749 => (0 => "11011110", 1 => "11000110", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            3750 => (0 => "11000110", 1 => "11001010", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            3751 => (0 => "11001010", 1 => "11001100", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            3752 => (0 => "11001100", 1 => "11001111", 2 => "11001110", 3 => "11001110", 4 => "11111111"),
            3753 => (0 => "01001111", 1 => "10001111", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            3754 => (0 => "10001111", 1 => "11101111", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            3755 => (0 => "11101111", 1 => "11011111", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            3756 => (0 => "11011111", 1 => "11000111", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            3757 => (0 => "11000111", 1 => "11001011", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            3758 => (0 => "11001011", 1 => "11001101", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            3759 => (0 => "11001101", 1 => "11001110", 2 => "11001111", 3 => "11001111", 4 => "11111111"),
            3760 => (0 => "01010000", 1 => "10010000", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            3761 => (0 => "10010000", 1 => "11110000", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            3762 => (0 => "11110000", 1 => "11000000", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            3763 => (0 => "11000000", 1 => "11011000", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            3764 => (0 => "11011000", 1 => "11010100", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            3765 => (0 => "11010100", 1 => "11010010", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            3766 => (0 => "11010010", 1 => "11010001", 2 => "11010000", 3 => "11010000", 4 => "11111111"),
            3767 => (0 => "01010001", 1 => "10010001", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            3768 => (0 => "10010001", 1 => "11110001", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            3769 => (0 => "11110001", 1 => "11000001", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            3770 => (0 => "11000001", 1 => "11011001", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            3771 => (0 => "11011001", 1 => "11010101", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            3772 => (0 => "11010101", 1 => "11010011", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            3773 => (0 => "11010011", 1 => "11010000", 2 => "11010001", 3 => "11010001", 4 => "11111111"),
            3774 => (0 => "01010010", 1 => "10010010", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            3775 => (0 => "10010010", 1 => "11110010", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            3776 => (0 => "11110010", 1 => "11000010", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            3777 => (0 => "11000010", 1 => "11011010", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            3778 => (0 => "11011010", 1 => "11010110", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            3779 => (0 => "11010110", 1 => "11010000", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            3780 => (0 => "11010000", 1 => "11010011", 2 => "11010010", 3 => "11010010", 4 => "11111111"),
            3781 => (0 => "01010011", 1 => "10010011", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            3782 => (0 => "10010011", 1 => "11110011", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            3783 => (0 => "11110011", 1 => "11000011", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            3784 => (0 => "11000011", 1 => "11011011", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            3785 => (0 => "11011011", 1 => "11010111", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            3786 => (0 => "11010111", 1 => "11010001", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            3787 => (0 => "11010001", 1 => "11010010", 2 => "11010011", 3 => "11010011", 4 => "11111111"),
            3788 => (0 => "01010100", 1 => "10010100", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            3789 => (0 => "10010100", 1 => "11110100", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            3790 => (0 => "11110100", 1 => "11000100", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            3791 => (0 => "11000100", 1 => "11011100", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            3792 => (0 => "11011100", 1 => "11010000", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            3793 => (0 => "11010000", 1 => "11010110", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            3794 => (0 => "11010110", 1 => "11010101", 2 => "11010100", 3 => "11010100", 4 => "11111111"),
            3795 => (0 => "01010101", 1 => "10010101", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            3796 => (0 => "10010101", 1 => "11110101", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            3797 => (0 => "11110101", 1 => "11000101", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            3798 => (0 => "11000101", 1 => "11011101", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            3799 => (0 => "11011101", 1 => "11010001", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            3800 => (0 => "11010001", 1 => "11010111", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            3801 => (0 => "11010111", 1 => "11010100", 2 => "11010101", 3 => "11010101", 4 => "11111111"),
            3802 => (0 => "01010110", 1 => "10010110", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            3803 => (0 => "10010110", 1 => "11110110", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            3804 => (0 => "11110110", 1 => "11000110", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            3805 => (0 => "11000110", 1 => "11011110", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            3806 => (0 => "11011110", 1 => "11010010", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            3807 => (0 => "11010010", 1 => "11010100", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            3808 => (0 => "11010100", 1 => "11010111", 2 => "11010110", 3 => "11010110", 4 => "11111111"),
            3809 => (0 => "01010111", 1 => "10010111", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            3810 => (0 => "10010111", 1 => "11110111", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            3811 => (0 => "11110111", 1 => "11000111", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            3812 => (0 => "11000111", 1 => "11011111", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            3813 => (0 => "11011111", 1 => "11010011", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            3814 => (0 => "11010011", 1 => "11010101", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            3815 => (0 => "11010101", 1 => "11010110", 2 => "11010111", 3 => "11010111", 4 => "11111111"),
            3816 => (0 => "01011000", 1 => "10011000", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            3817 => (0 => "10011000", 1 => "11111000", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            3818 => (0 => "11111000", 1 => "11001000", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            3819 => (0 => "11001000", 1 => "11010000", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            3820 => (0 => "11010000", 1 => "11011100", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            3821 => (0 => "11011100", 1 => "11011010", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            3822 => (0 => "11011010", 1 => "11011001", 2 => "11011000", 3 => "11011000", 4 => "11111111"),
            3823 => (0 => "01011001", 1 => "10011001", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            3824 => (0 => "10011001", 1 => "11111001", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            3825 => (0 => "11111001", 1 => "11001001", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            3826 => (0 => "11001001", 1 => "11010001", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            3827 => (0 => "11010001", 1 => "11011101", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            3828 => (0 => "11011101", 1 => "11011011", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            3829 => (0 => "11011011", 1 => "11011000", 2 => "11011001", 3 => "11011001", 4 => "11111111"),
            3830 => (0 => "01011010", 1 => "10011010", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            3831 => (0 => "10011010", 1 => "11111010", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            3832 => (0 => "11111010", 1 => "11001010", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            3833 => (0 => "11001010", 1 => "11010010", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            3834 => (0 => "11010010", 1 => "11011110", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            3835 => (0 => "11011110", 1 => "11011000", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            3836 => (0 => "11011000", 1 => "11011011", 2 => "11011010", 3 => "11011010", 4 => "11111111"),
            3837 => (0 => "01011011", 1 => "10011011", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            3838 => (0 => "10011011", 1 => "11111011", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            3839 => (0 => "11111011", 1 => "11001011", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            3840 => (0 => "11001011", 1 => "11010011", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            3841 => (0 => "11010011", 1 => "11011111", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            3842 => (0 => "11011111", 1 => "11011001", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            3843 => (0 => "11011001", 1 => "11011010", 2 => "11011011", 3 => "11011011", 4 => "11111111"),
            3844 => (0 => "01011100", 1 => "10011100", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            3845 => (0 => "10011100", 1 => "11111100", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            3846 => (0 => "11111100", 1 => "11001100", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            3847 => (0 => "11001100", 1 => "11010100", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            3848 => (0 => "11010100", 1 => "11011000", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            3849 => (0 => "11011000", 1 => "11011110", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            3850 => (0 => "11011110", 1 => "11011101", 2 => "11011100", 3 => "11011100", 4 => "11111111"),
            3851 => (0 => "01011101", 1 => "10011101", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            3852 => (0 => "10011101", 1 => "11111101", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            3853 => (0 => "11111101", 1 => "11001101", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            3854 => (0 => "11001101", 1 => "11010101", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            3855 => (0 => "11010101", 1 => "11011001", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            3856 => (0 => "11011001", 1 => "11011111", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            3857 => (0 => "11011111", 1 => "11011100", 2 => "11011101", 3 => "11011101", 4 => "11111111"),
            3858 => (0 => "01011110", 1 => "10011110", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            3859 => (0 => "10011110", 1 => "11111110", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            3860 => (0 => "11111110", 1 => "11001110", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            3861 => (0 => "11001110", 1 => "11010110", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            3862 => (0 => "11010110", 1 => "11011010", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            3863 => (0 => "11011010", 1 => "11011100", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            3864 => (0 => "11011100", 1 => "11011111", 2 => "11011110", 3 => "11011110", 4 => "11111111"),
            3865 => (0 => "01011111", 1 => "10011111", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            3866 => (0 => "10011111", 1 => "11111111", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            3867 => (0 => "11111111", 1 => "11001111", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            3868 => (0 => "11001111", 1 => "11010111", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            3869 => (0 => "11010111", 1 => "11011011", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            3870 => (0 => "11011011", 1 => "11011101", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            3871 => (0 => "11011101", 1 => "11011110", 2 => "11011111", 3 => "11011111", 4 => "11111111"),
            3872 => (0 => "01100000", 1 => "10100000", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            3873 => (0 => "10100000", 1 => "11000000", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            3874 => (0 => "11000000", 1 => "11110000", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            3875 => (0 => "11110000", 1 => "11101000", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            3876 => (0 => "11101000", 1 => "11100100", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            3877 => (0 => "11100100", 1 => "11100010", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            3878 => (0 => "11100010", 1 => "11100001", 2 => "11100000", 3 => "11100000", 4 => "11111111"),
            3879 => (0 => "01100001", 1 => "10100001", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            3880 => (0 => "10100001", 1 => "11000001", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            3881 => (0 => "11000001", 1 => "11110001", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            3882 => (0 => "11110001", 1 => "11101001", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            3883 => (0 => "11101001", 1 => "11100101", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            3884 => (0 => "11100101", 1 => "11100011", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            3885 => (0 => "11100011", 1 => "11100000", 2 => "11100001", 3 => "11100001", 4 => "11111111"),
            3886 => (0 => "01100010", 1 => "10100010", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            3887 => (0 => "10100010", 1 => "11000010", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            3888 => (0 => "11000010", 1 => "11110010", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            3889 => (0 => "11110010", 1 => "11101010", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            3890 => (0 => "11101010", 1 => "11100110", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            3891 => (0 => "11100110", 1 => "11100000", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            3892 => (0 => "11100000", 1 => "11100011", 2 => "11100010", 3 => "11100010", 4 => "11111111"),
            3893 => (0 => "01100011", 1 => "10100011", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            3894 => (0 => "10100011", 1 => "11000011", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            3895 => (0 => "11000011", 1 => "11110011", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            3896 => (0 => "11110011", 1 => "11101011", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            3897 => (0 => "11101011", 1 => "11100111", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            3898 => (0 => "11100111", 1 => "11100001", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            3899 => (0 => "11100001", 1 => "11100010", 2 => "11100011", 3 => "11100011", 4 => "11111111"),
            3900 => (0 => "01100100", 1 => "10100100", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            3901 => (0 => "10100100", 1 => "11000100", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            3902 => (0 => "11000100", 1 => "11110100", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            3903 => (0 => "11110100", 1 => "11101100", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            3904 => (0 => "11101100", 1 => "11100000", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            3905 => (0 => "11100000", 1 => "11100110", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            3906 => (0 => "11100110", 1 => "11100101", 2 => "11100100", 3 => "11100100", 4 => "11111111"),
            3907 => (0 => "01100101", 1 => "10100101", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            3908 => (0 => "10100101", 1 => "11000101", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            3909 => (0 => "11000101", 1 => "11110101", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            3910 => (0 => "11110101", 1 => "11101101", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            3911 => (0 => "11101101", 1 => "11100001", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            3912 => (0 => "11100001", 1 => "11100111", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            3913 => (0 => "11100111", 1 => "11100100", 2 => "11100101", 3 => "11100101", 4 => "11111111"),
            3914 => (0 => "01100110", 1 => "10100110", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            3915 => (0 => "10100110", 1 => "11000110", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            3916 => (0 => "11000110", 1 => "11110110", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            3917 => (0 => "11110110", 1 => "11101110", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            3918 => (0 => "11101110", 1 => "11100010", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            3919 => (0 => "11100010", 1 => "11100100", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            3920 => (0 => "11100100", 1 => "11100111", 2 => "11100110", 3 => "11100110", 4 => "11111111"),
            3921 => (0 => "01100111", 1 => "10100111", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            3922 => (0 => "10100111", 1 => "11000111", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            3923 => (0 => "11000111", 1 => "11110111", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            3924 => (0 => "11110111", 1 => "11101111", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            3925 => (0 => "11101111", 1 => "11100011", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            3926 => (0 => "11100011", 1 => "11100101", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            3927 => (0 => "11100101", 1 => "11100110", 2 => "11100111", 3 => "11100111", 4 => "11111111"),
            3928 => (0 => "01101000", 1 => "10101000", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            3929 => (0 => "10101000", 1 => "11001000", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            3930 => (0 => "11001000", 1 => "11111000", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            3931 => (0 => "11111000", 1 => "11100000", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            3932 => (0 => "11100000", 1 => "11101100", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            3933 => (0 => "11101100", 1 => "11101010", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            3934 => (0 => "11101010", 1 => "11101001", 2 => "11101000", 3 => "11101000", 4 => "11111111"),
            3935 => (0 => "01101001", 1 => "10101001", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            3936 => (0 => "10101001", 1 => "11001001", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            3937 => (0 => "11001001", 1 => "11111001", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            3938 => (0 => "11111001", 1 => "11100001", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            3939 => (0 => "11100001", 1 => "11101101", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            3940 => (0 => "11101101", 1 => "11101011", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            3941 => (0 => "11101011", 1 => "11101000", 2 => "11101001", 3 => "11101001", 4 => "11111111"),
            3942 => (0 => "01101010", 1 => "10101010", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            3943 => (0 => "10101010", 1 => "11001010", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            3944 => (0 => "11001010", 1 => "11111010", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            3945 => (0 => "11111010", 1 => "11100010", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            3946 => (0 => "11100010", 1 => "11101110", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            3947 => (0 => "11101110", 1 => "11101000", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            3948 => (0 => "11101000", 1 => "11101011", 2 => "11101010", 3 => "11101010", 4 => "11111111"),
            3949 => (0 => "01101011", 1 => "10101011", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            3950 => (0 => "10101011", 1 => "11001011", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            3951 => (0 => "11001011", 1 => "11111011", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            3952 => (0 => "11111011", 1 => "11100011", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            3953 => (0 => "11100011", 1 => "11101111", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            3954 => (0 => "11101111", 1 => "11101001", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            3955 => (0 => "11101001", 1 => "11101010", 2 => "11101011", 3 => "11101011", 4 => "11111111"),
            3956 => (0 => "01101100", 1 => "10101100", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            3957 => (0 => "10101100", 1 => "11001100", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            3958 => (0 => "11001100", 1 => "11111100", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            3959 => (0 => "11111100", 1 => "11100100", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            3960 => (0 => "11100100", 1 => "11101000", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            3961 => (0 => "11101000", 1 => "11101110", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            3962 => (0 => "11101110", 1 => "11101101", 2 => "11101100", 3 => "11101100", 4 => "11111111"),
            3963 => (0 => "01101101", 1 => "10101101", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            3964 => (0 => "10101101", 1 => "11001101", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            3965 => (0 => "11001101", 1 => "11111101", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            3966 => (0 => "11111101", 1 => "11100101", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            3967 => (0 => "11100101", 1 => "11101001", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            3968 => (0 => "11101001", 1 => "11101111", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            3969 => (0 => "11101111", 1 => "11101100", 2 => "11101101", 3 => "11101101", 4 => "11111111"),
            3970 => (0 => "01101110", 1 => "10101110", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            3971 => (0 => "10101110", 1 => "11001110", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            3972 => (0 => "11001110", 1 => "11111110", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            3973 => (0 => "11111110", 1 => "11100110", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            3974 => (0 => "11100110", 1 => "11101010", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            3975 => (0 => "11101010", 1 => "11101100", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            3976 => (0 => "11101100", 1 => "11101111", 2 => "11101110", 3 => "11101110", 4 => "11111111"),
            3977 => (0 => "01101111", 1 => "10101111", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            3978 => (0 => "10101111", 1 => "11001111", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            3979 => (0 => "11001111", 1 => "11111111", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            3980 => (0 => "11111111", 1 => "11100111", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            3981 => (0 => "11100111", 1 => "11101011", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            3982 => (0 => "11101011", 1 => "11101101", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            3983 => (0 => "11101101", 1 => "11101110", 2 => "11101111", 3 => "11101111", 4 => "11111111"),
            3984 => (0 => "01110000", 1 => "10110000", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            3985 => (0 => "10110000", 1 => "11010000", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            3986 => (0 => "11010000", 1 => "11100000", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            3987 => (0 => "11100000", 1 => "11111000", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            3988 => (0 => "11111000", 1 => "11110100", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            3989 => (0 => "11110100", 1 => "11110010", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            3990 => (0 => "11110010", 1 => "11110001", 2 => "11110000", 3 => "11110000", 4 => "11111111"),
            3991 => (0 => "01110001", 1 => "10110001", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            3992 => (0 => "10110001", 1 => "11010001", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            3993 => (0 => "11010001", 1 => "11100001", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            3994 => (0 => "11100001", 1 => "11111001", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            3995 => (0 => "11111001", 1 => "11110101", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            3996 => (0 => "11110101", 1 => "11110011", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            3997 => (0 => "11110011", 1 => "11110000", 2 => "11110001", 3 => "11110001", 4 => "11111111"),
            3998 => (0 => "01110010", 1 => "10110010", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            3999 => (0 => "10110010", 1 => "11010010", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            4000 => (0 => "11010010", 1 => "11100010", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            4001 => (0 => "11100010", 1 => "11111010", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            4002 => (0 => "11111010", 1 => "11110110", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            4003 => (0 => "11110110", 1 => "11110000", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            4004 => (0 => "11110000", 1 => "11110011", 2 => "11110010", 3 => "11110010", 4 => "11111111"),
            4005 => (0 => "01110011", 1 => "10110011", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            4006 => (0 => "10110011", 1 => "11010011", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            4007 => (0 => "11010011", 1 => "11100011", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            4008 => (0 => "11100011", 1 => "11111011", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            4009 => (0 => "11111011", 1 => "11110111", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            4010 => (0 => "11110111", 1 => "11110001", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            4011 => (0 => "11110001", 1 => "11110010", 2 => "11110011", 3 => "11110011", 4 => "11111111"),
            4012 => (0 => "01110100", 1 => "10110100", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            4013 => (0 => "10110100", 1 => "11010100", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            4014 => (0 => "11010100", 1 => "11100100", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            4015 => (0 => "11100100", 1 => "11111100", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            4016 => (0 => "11111100", 1 => "11110000", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            4017 => (0 => "11110000", 1 => "11110110", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            4018 => (0 => "11110110", 1 => "11110101", 2 => "11110100", 3 => "11110100", 4 => "11111111"),
            4019 => (0 => "01110101", 1 => "10110101", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            4020 => (0 => "10110101", 1 => "11010101", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            4021 => (0 => "11010101", 1 => "11100101", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            4022 => (0 => "11100101", 1 => "11111101", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            4023 => (0 => "11111101", 1 => "11110001", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            4024 => (0 => "11110001", 1 => "11110111", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            4025 => (0 => "11110111", 1 => "11110100", 2 => "11110101", 3 => "11110101", 4 => "11111111"),
            4026 => (0 => "01110110", 1 => "10110110", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            4027 => (0 => "10110110", 1 => "11010110", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            4028 => (0 => "11010110", 1 => "11100110", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            4029 => (0 => "11100110", 1 => "11111110", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            4030 => (0 => "11111110", 1 => "11110010", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            4031 => (0 => "11110010", 1 => "11110100", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            4032 => (0 => "11110100", 1 => "11110111", 2 => "11110110", 3 => "11110110", 4 => "11111111"),
            4033 => (0 => "01110111", 1 => "10110111", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            4034 => (0 => "10110111", 1 => "11010111", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            4035 => (0 => "11010111", 1 => "11100111", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            4036 => (0 => "11100111", 1 => "11111111", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            4037 => (0 => "11111111", 1 => "11110011", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            4038 => (0 => "11110011", 1 => "11110101", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            4039 => (0 => "11110101", 1 => "11110110", 2 => "11110111", 3 => "11110111", 4 => "11111111"),
            4040 => (0 => "01111000", 1 => "10111000", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            4041 => (0 => "10111000", 1 => "11011000", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            4042 => (0 => "11011000", 1 => "11101000", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            4043 => (0 => "11101000", 1 => "11110000", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            4044 => (0 => "11110000", 1 => "11111100", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            4045 => (0 => "11111100", 1 => "11111010", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            4046 => (0 => "11111010", 1 => "11111001", 2 => "11111000", 3 => "11111000", 4 => "11111111"),
            4047 => (0 => "01111001", 1 => "10111001", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            4048 => (0 => "10111001", 1 => "11011001", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            4049 => (0 => "11011001", 1 => "11101001", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            4050 => (0 => "11101001", 1 => "11110001", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            4051 => (0 => "11110001", 1 => "11111101", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            4052 => (0 => "11111101", 1 => "11111011", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            4053 => (0 => "11111011", 1 => "11111000", 2 => "11111001", 3 => "11111001", 4 => "11111111"),
            4054 => (0 => "01111010", 1 => "10111010", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            4055 => (0 => "10111010", 1 => "11011010", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            4056 => (0 => "11011010", 1 => "11101010", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            4057 => (0 => "11101010", 1 => "11110010", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            4058 => (0 => "11110010", 1 => "11111110", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            4059 => (0 => "11111110", 1 => "11111000", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            4060 => (0 => "11111000", 1 => "11111011", 2 => "11111010", 3 => "11111010", 4 => "11111111"),
            4061 => (0 => "01111011", 1 => "10111011", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            4062 => (0 => "10111011", 1 => "11011011", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            4063 => (0 => "11011011", 1 => "11101011", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            4064 => (0 => "11101011", 1 => "11110011", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            4065 => (0 => "11110011", 1 => "11111111", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            4066 => (0 => "11111111", 1 => "11111001", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            4067 => (0 => "11111001", 1 => "11111010", 2 => "11111011", 3 => "11111011", 4 => "11111111"),
            4068 => (0 => "01111100", 1 => "10111100", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            4069 => (0 => "10111100", 1 => "11011100", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            4070 => (0 => "11011100", 1 => "11101100", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            4071 => (0 => "11101100", 1 => "11110100", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            4072 => (0 => "11110100", 1 => "11111000", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            4073 => (0 => "11111000", 1 => "11111110", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            4074 => (0 => "11111110", 1 => "11111101", 2 => "11111100", 3 => "11111100", 4 => "11111111"),
            4075 => (0 => "01111101", 1 => "10111101", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            4076 => (0 => "10111101", 1 => "11011101", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            4077 => (0 => "11011101", 1 => "11101101", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            4078 => (0 => "11101101", 1 => "11110101", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            4079 => (0 => "11110101", 1 => "11111001", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            4080 => (0 => "11111001", 1 => "11111111", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            4081 => (0 => "11111111", 1 => "11111100", 2 => "11111101", 3 => "11111101", 4 => "11111111"),
            4082 => (0 => "01111110", 1 => "10111110", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            4083 => (0 => "10111110", 1 => "11011110", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            4084 => (0 => "11011110", 1 => "11101110", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            4085 => (0 => "11101110", 1 => "11110110", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            4086 => (0 => "11110110", 1 => "11111010", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            4087 => (0 => "11111010", 1 => "11111100", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            4088 => (0 => "11111100", 1 => "11111111", 2 => "11111110", 3 => "11111110", 4 => "11111111"),
            4089 => (0 => "01111111", 1 => "10111111", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            4090 => (0 => "10111111", 1 => "11011111", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            4091 => (0 => "11011111", 1 => "11101111", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            4092 => (0 => "11101111", 1 => "11110111", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            4093 => (0 => "11110111", 1 => "11111011", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            4094 => (0 => "11111011", 1 => "11111101", 2 => "11111111", 3 => "11111111", 4 => "11111111"),
            4095 => (0 => "11111101", 1 => "11111110", 2 => "11111111", 3 => "11111111", 4 => "11111111")
    );
	
	-- 0 => "00000000" & "000"  & "0000",
	constant output : outputvect_t := (
	                0 => "000000000000000",
            1 => "000000010000111",
            2 => "000000100001001",
            3 => "000000110001110",
            4 => "000001000001010",
            5 => "000001010001101",
            6 => "000001100000011",
            7 => "000001110000100",
            8 => "000010000001011",
            9 => "000010010001100",
            10 => "000010100000010",
            11 => "000010110000101",
            12 => "000011000000001",
            13 => "000011010000110",
            14 => "000011100001000",
            15 => "000011110001111",
            16 => "000100000001100",
            17 => "000100010001011",
            18 => "000100100000101",
            19 => "000100110000010",
            20 => "000101000000110",
            21 => "000101010000001",
            22 => "000101100001111",
            23 => "000101110001000",
            24 => "000110000000111",
            25 => "000110010000000",
            26 => "000110100001110",
            27 => "000110110001001",
            28 => "000111000001101",
            29 => "000111010001010",
            30 => "000111100000100",
            31 => "000111110000011",
            32 => "001000000001101",
            33 => "001000010001010",
            34 => "001000100000100",
            35 => "001000110000011",
            36 => "001001000000111",
            37 => "001001010000000",
            38 => "001001100001110",
            39 => "001001110001001",
            40 => "001010000000110",
            41 => "001010010000001",
            42 => "001010100001111",
            43 => "001010110001000",
            44 => "001011000001100",
            45 => "001011010001011",
            46 => "001011100000101",
            47 => "001011110000010",
            48 => "001100000000001",
            49 => "001100010000110",
            50 => "001100100001000",
            51 => "001100110001111",
            52 => "001101000001011",
            53 => "001101010001100",
            54 => "001101100000010",
            55 => "001101110000101",
            56 => "001110000001010",
            57 => "001110010001101",
            58 => "001110100000011",
            59 => "001110110000100",
            60 => "001111000000000",
            61 => "001111010000111",
            62 => "001111100001001",
            63 => "001111110001110",
            64 => "010000000001110",
            65 => "010000010001001",
            66 => "010000100000111",
            67 => "010000110000000",
            68 => "010001000000100",
            69 => "010001010000011",
            70 => "010001100001101",
            71 => "010001110001010",
            72 => "010010000000101",
            73 => "010010010000010",
            74 => "010010100001100",
            75 => "010010110001011",
            76 => "010011000001111",
            77 => "010011010001000",
            78 => "010011100000110",
            79 => "010011110000001",
            80 => "010100000000010",
            81 => "010100010000101",
            82 => "010100100001011",
            83 => "010100110001100",
            84 => "010101000001000",
            85 => "010101010001111",
            86 => "010101100000001",
            87 => "010101110000110",
            88 => "010110000001001",
            89 => "010110010001110",
            90 => "010110100000000",
            91 => "010110110000111",
            92 => "010111000000011",
            93 => "010111010000100",
            94 => "010111100001010",
            95 => "010111110001101",
            96 => "011000000000011",
            97 => "011000010000100",
            98 => "011000100001010",
            99 => "011000110001101",
            100 => "011001000001001",
            101 => "011001010001110",
            102 => "011001100000000",
            103 => "011001110000111",
            104 => "011010000001000",
            105 => "011010010001111",
            106 => "011010100000001",
            107 => "011010110000110",
            108 => "011011000000010",
            109 => "011011010000101",
            110 => "011011100001011",
            111 => "011011110001100",
            112 => "011100000001111",
            113 => "011100010001000",
            114 => "011100100000110",
            115 => "011100110000001",
            116 => "011101000000101",
            117 => "011101010000010",
            118 => "011101100001100",
            119 => "011101110001011",
            120 => "011110000000100",
            121 => "011110010000011",
            122 => "011110100001101",
            123 => "011110110001010",
            124 => "011111000001110",
            125 => "011111010001001",
            126 => "011111100000111",
            127 => "011111110000000",
            128 => "100000000001111",
            129 => "100000010001000",
            130 => "100000100000110",
            131 => "100000110000001",
            132 => "100001000000101",
            133 => "100001010000010",
            134 => "100001100001100",
            135 => "100001110001011",
            136 => "100010000000100",
            137 => "100010010000011",
            138 => "100010100001101",
            139 => "100010110001010",
            140 => "100011000001110",
            141 => "100011010001001",
            142 => "100011100000111",
            143 => "100011110000000",
            144 => "100100000000011",
            145 => "100100010000100",
            146 => "100100100001010",
            147 => "100100110001101",
            148 => "100101000001001",
            149 => "100101010001110",
            150 => "100101100000000",
            151 => "100101110000111",
            152 => "100110000001000",
            153 => "100110010001111",
            154 => "100110100000001",
            155 => "100110110000110",
            156 => "100111000000010",
            157 => "100111010000101",
            158 => "100111100001011",
            159 => "100111110001100",
            160 => "101000000000010",
            161 => "101000010000101",
            162 => "101000100001011",
            163 => "101000110001100",
            164 => "101001000001000",
            165 => "101001010001111",
            166 => "101001100000001",
            167 => "101001110000110",
            168 => "101010000001001",
            169 => "101010010001110",
            170 => "101010100000000",
            171 => "101010110000111",
            172 => "101011000000011",
            173 => "101011010000100",
            174 => "101011100001010",
            175 => "101011110001101",
            176 => "101100000001110",
            177 => "101100010001001",
            178 => "101100100000111",
            179 => "101100110000000",
            180 => "101101000000100",
            181 => "101101010000011",
            182 => "101101100001101",
            183 => "101101110001010",
            184 => "101110000000101",
            185 => "101110010000010",
            186 => "101110100001100",
            187 => "101110110001011",
            188 => "101111000001111",
            189 => "101111010001000",
            190 => "101111100000110",
            191 => "101111110000001",
            192 => "110000000000001",
            193 => "110000010000110",
            194 => "110000100001000",
            195 => "110000110001111",
            196 => "110001000001011",
            197 => "110001010001100",
            198 => "110001100000010",
            199 => "110001110000101",
            200 => "110010000001010",
            201 => "110010010001101",
            202 => "110010100000011",
            203 => "110010110000100",
            204 => "110011000000000",
            205 => "110011010000111",
            206 => "110011100001001",
            207 => "110011110001110",
            208 => "110100000001101",
            209 => "110100010001010",
            210 => "110100100000100",
            211 => "110100110000011",
            212 => "110101000000111",
            213 => "110101010000000",
            214 => "110101100001110",
            215 => "110101110001001",
            216 => "110110000000110",
            217 => "110110010000001",
            218 => "110110100001111",
            219 => "110110110001000",
            220 => "110111000001100",
            221 => "110111010001011",
            222 => "110111100000101",
            223 => "110111110000010",
            224 => "111000000001100",
            225 => "111000010001011",
            226 => "111000100000101",
            227 => "111000110000010",
            228 => "111001000000110",
            229 => "111001010000001",
            230 => "111001100001111",
            231 => "111001110001000",
            232 => "111010000000111",
            233 => "111010010000000",
            234 => "111010100001110",
            235 => "111010110001001",
            236 => "111011000001101",
            237 => "111011010001010",
            238 => "111011100000100",
            239 => "111011110000011",
            240 => "111100000000000",
            241 => "111100010000111",
            242 => "111100100001001",
            243 => "111100110001110",
            244 => "111101000001010",
            245 => "111101010001101",
            246 => "111101100000011",
            247 => "111101110000100",
            248 => "111110000001011",
            249 => "111110010001100",
            250 => "111110100000010",
            251 => "111110110000101",
            252 => "111111000000001",
            253 => "111111010000110",
            254 => "111111100001000",
            255 => "111111110001111",
            256 => "000000000010011",
            257 => "000000000010011",
            258 => "000000000010011",
            259 => "000000000010011",
            260 => "000000000010011",
            261 => "000000000010011",
            262 => "000000000010011",
            263 => "000000000010011",
            264 => "000000010010100",
            265 => "000000010010100",
            266 => "000000010010100",
            267 => "000000010010100",
            268 => "000000010010100",
            269 => "000000010010100",
            270 => "000000010010100",
            271 => "000000010010100",
            272 => "000000100011010",
            273 => "000000100011010",
            274 => "000000100011010",
            275 => "000000100011010",
            276 => "000000100011010",
            277 => "000000100011010",
            278 => "000000100011010",
            279 => "000000100011010",
            280 => "000000110011101",
            281 => "000000110011101",
            282 => "000000110011101",
            283 => "000000110011101",
            284 => "000000110011101",
            285 => "000000110011101",
            286 => "000000110011101",
            287 => "000000110011101",
            288 => "000001000011001",
            289 => "000001000011001",
            290 => "000001000011001",
            291 => "000001000011001",
            292 => "000001000011001",
            293 => "000001000011001",
            294 => "000001000011001",
            295 => "000001000011001",
            296 => "000001010011110",
            297 => "000001010011110",
            298 => "000001010011110",
            299 => "000001010011110",
            300 => "000001010011110",
            301 => "000001010011110",
            302 => "000001010011110",
            303 => "000001010011110",
            304 => "000001100010000",
            305 => "000001100010000",
            306 => "000001100010000",
            307 => "000001100010000",
            308 => "000001100010000",
            309 => "000001100010000",
            310 => "000001100010000",
            311 => "000001100010000",
            312 => "000001110010111",
            313 => "000001110010111",
            314 => "000001110010111",
            315 => "000001110010111",
            316 => "000001110010111",
            317 => "000001110010111",
            318 => "000001110010111",
            319 => "000001110010111",
            320 => "000010000011000",
            321 => "000010000011000",
            322 => "000010000011000",
            323 => "000010000011000",
            324 => "000010000011000",
            325 => "000010000011000",
            326 => "000010000011000",
            327 => "000010000011000",
            328 => "000010010011111",
            329 => "000010010011111",
            330 => "000010010011111",
            331 => "000010010011111",
            332 => "000010010011111",
            333 => "000010010011111",
            334 => "000010010011111",
            335 => "000010010011111",
            336 => "000010100010001",
            337 => "000010100010001",
            338 => "000010100010001",
            339 => "000010100010001",
            340 => "000010100010001",
            341 => "000010100010001",
            342 => "000010100010001",
            343 => "000010100010001",
            344 => "000010110010110",
            345 => "000010110010110",
            346 => "000010110010110",
            347 => "000010110010110",
            348 => "000010110010110",
            349 => "000010110010110",
            350 => "000010110010110",
            351 => "000010110010110",
            352 => "000011000010010",
            353 => "000011000010010",
            354 => "000011000010010",
            355 => "000011000010010",
            356 => "000011000010010",
            357 => "000011000010010",
            358 => "000011000010010",
            359 => "000011000010010",
            360 => "000011010010101",
            361 => "000011010010101",
            362 => "000011010010101",
            363 => "000011010010101",
            364 => "000011010010101",
            365 => "000011010010101",
            366 => "000011010010101",
            367 => "000011010010101",
            368 => "000011100011011",
            369 => "000011100011011",
            370 => "000011100011011",
            371 => "000011100011011",
            372 => "000011100011011",
            373 => "000011100011011",
            374 => "000011100011011",
            375 => "000011100011011",
            376 => "000011110011100",
            377 => "000011110011100",
            378 => "000011110011100",
            379 => "000011110011100",
            380 => "000011110011100",
            381 => "000011110011100",
            382 => "000011110011100",
            383 => "000011110011100",
            384 => "000100000011111",
            385 => "000100000011111",
            386 => "000100000011111",
            387 => "000100000011111",
            388 => "000100000011111",
            389 => "000100000011111",
            390 => "000100000011111",
            391 => "000100000011111",
            392 => "000100010011000",
            393 => "000100010011000",
            394 => "000100010011000",
            395 => "000100010011000",
            396 => "000100010011000",
            397 => "000100010011000",
            398 => "000100010011000",
            399 => "000100010011000",
            400 => "000100100010110",
            401 => "000100100010110",
            402 => "000100100010110",
            403 => "000100100010110",
            404 => "000100100010110",
            405 => "000100100010110",
            406 => "000100100010110",
            407 => "000100100010110",
            408 => "000100110010001",
            409 => "000100110010001",
            410 => "000100110010001",
            411 => "000100110010001",
            412 => "000100110010001",
            413 => "000100110010001",
            414 => "000100110010001",
            415 => "000100110010001",
            416 => "000101000010101",
            417 => "000101000010101",
            418 => "000101000010101",
            419 => "000101000010101",
            420 => "000101000010101",
            421 => "000101000010101",
            422 => "000101000010101",
            423 => "000101000010101",
            424 => "000101010010010",
            425 => "000101010010010",
            426 => "000101010010010",
            427 => "000101010010010",
            428 => "000101010010010",
            429 => "000101010010010",
            430 => "000101010010010",
            431 => "000101010010010",
            432 => "000101100011100",
            433 => "000101100011100",
            434 => "000101100011100",
            435 => "000101100011100",
            436 => "000101100011100",
            437 => "000101100011100",
            438 => "000101100011100",
            439 => "000101100011100",
            440 => "000101110011011",
            441 => "000101110011011",
            442 => "000101110011011",
            443 => "000101110011011",
            444 => "000101110011011",
            445 => "000101110011011",
            446 => "000101110011011",
            447 => "000101110011011",
            448 => "000110000010100",
            449 => "000110000010100",
            450 => "000110000010100",
            451 => "000110000010100",
            452 => "000110000010100",
            453 => "000110000010100",
            454 => "000110000010100",
            455 => "000110000010100",
            456 => "000110010010011",
            457 => "000110010010011",
            458 => "000110010010011",
            459 => "000110010010011",
            460 => "000110010010011",
            461 => "000110010010011",
            462 => "000110010010011",
            463 => "000110010010011",
            464 => "000110100011101",
            465 => "000110100011101",
            466 => "000110100011101",
            467 => "000110100011101",
            468 => "000110100011101",
            469 => "000110100011101",
            470 => "000110100011101",
            471 => "000110100011101",
            472 => "000110110011010",
            473 => "000110110011010",
            474 => "000110110011010",
            475 => "000110110011010",
            476 => "000110110011010",
            477 => "000110110011010",
            478 => "000110110011010",
            479 => "000110110011010",
            480 => "000111000011110",
            481 => "000111000011110",
            482 => "000111000011110",
            483 => "000111000011110",
            484 => "000111000011110",
            485 => "000111000011110",
            486 => "000111000011110",
            487 => "000111000011110",
            488 => "000111010011001",
            489 => "000111010011001",
            490 => "000111010011001",
            491 => "000111010011001",
            492 => "000111010011001",
            493 => "000111010011001",
            494 => "000111010011001",
            495 => "000111010011001",
            496 => "000111100010111",
            497 => "000111100010111",
            498 => "000111100010111",
            499 => "000111100010111",
            500 => "000111100010111",
            501 => "000111100010111",
            502 => "000111100010111",
            503 => "000111100010111",
            504 => "000111110010000",
            505 => "000111110010000",
            506 => "000111110010000",
            507 => "000111110010000",
            508 => "000111110010000",
            509 => "000111110010000",
            510 => "000111110010000",
            511 => "000111110010000",
            512 => "001000000011110",
            513 => "001000000011110",
            514 => "001000000011110",
            515 => "001000000011110",
            516 => "001000000011110",
            517 => "001000000011110",
            518 => "001000000011110",
            519 => "001000000011110",
            520 => "001000010011001",
            521 => "001000010011001",
            522 => "001000010011001",
            523 => "001000010011001",
            524 => "001000010011001",
            525 => "001000010011001",
            526 => "001000010011001",
            527 => "001000010011001",
            528 => "001000100010111",
            529 => "001000100010111",
            530 => "001000100010111",
            531 => "001000100010111",
            532 => "001000100010111",
            533 => "001000100010111",
            534 => "001000100010111",
            535 => "001000100010111",
            536 => "001000110010000",
            537 => "001000110010000",
            538 => "001000110010000",
            539 => "001000110010000",
            540 => "001000110010000",
            541 => "001000110010000",
            542 => "001000110010000",
            543 => "001000110010000",
            544 => "001001000010100",
            545 => "001001000010100",
            546 => "001001000010100",
            547 => "001001000010100",
            548 => "001001000010100",
            549 => "001001000010100",
            550 => "001001000010100",
            551 => "001001000010100",
            552 => "001001010010011",
            553 => "001001010010011",
            554 => "001001010010011",
            555 => "001001010010011",
            556 => "001001010010011",
            557 => "001001010010011",
            558 => "001001010010011",
            559 => "001001010010011",
            560 => "001001100011101",
            561 => "001001100011101",
            562 => "001001100011101",
            563 => "001001100011101",
            564 => "001001100011101",
            565 => "001001100011101",
            566 => "001001100011101",
            567 => "001001100011101",
            568 => "001001110011010",
            569 => "001001110011010",
            570 => "001001110011010",
            571 => "001001110011010",
            572 => "001001110011010",
            573 => "001001110011010",
            574 => "001001110011010",
            575 => "001001110011010",
            576 => "001010000010101",
            577 => "001010000010101",
            578 => "001010000010101",
            579 => "001010000010101",
            580 => "001010000010101",
            581 => "001010000010101",
            582 => "001010000010101",
            583 => "001010000010101",
            584 => "001010010010010",
            585 => "001010010010010",
            586 => "001010010010010",
            587 => "001010010010010",
            588 => "001010010010010",
            589 => "001010010010010",
            590 => "001010010010010",
            591 => "001010010010010",
            592 => "001010100011100",
            593 => "001010100011100",
            594 => "001010100011100",
            595 => "001010100011100",
            596 => "001010100011100",
            597 => "001010100011100",
            598 => "001010100011100",
            599 => "001010100011100",
            600 => "001010110011011",
            601 => "001010110011011",
            602 => "001010110011011",
            603 => "001010110011011",
            604 => "001010110011011",
            605 => "001010110011011",
            606 => "001010110011011",
            607 => "001010110011011",
            608 => "001011000011111",
            609 => "001011000011111",
            610 => "001011000011111",
            611 => "001011000011111",
            612 => "001011000011111",
            613 => "001011000011111",
            614 => "001011000011111",
            615 => "001011000011111",
            616 => "001011010011000",
            617 => "001011010011000",
            618 => "001011010011000",
            619 => "001011010011000",
            620 => "001011010011000",
            621 => "001011010011000",
            622 => "001011010011000",
            623 => "001011010011000",
            624 => "001011100010110",
            625 => "001011100010110",
            626 => "001011100010110",
            627 => "001011100010110",
            628 => "001011100010110",
            629 => "001011100010110",
            630 => "001011100010110",
            631 => "001011100010110",
            632 => "001011110010001",
            633 => "001011110010001",
            634 => "001011110010001",
            635 => "001011110010001",
            636 => "001011110010001",
            637 => "001011110010001",
            638 => "001011110010001",
            639 => "001011110010001",
            640 => "001100000010010",
            641 => "001100000010010",
            642 => "001100000010010",
            643 => "001100000010010",
            644 => "001100000010010",
            645 => "001100000010010",
            646 => "001100000010010",
            647 => "001100000010010",
            648 => "001100010010101",
            649 => "001100010010101",
            650 => "001100010010101",
            651 => "001100010010101",
            652 => "001100010010101",
            653 => "001100010010101",
            654 => "001100010010101",
            655 => "001100010010101",
            656 => "001100100011011",
            657 => "001100100011011",
            658 => "001100100011011",
            659 => "001100100011011",
            660 => "001100100011011",
            661 => "001100100011011",
            662 => "001100100011011",
            663 => "001100100011011",
            664 => "001100110011100",
            665 => "001100110011100",
            666 => "001100110011100",
            667 => "001100110011100",
            668 => "001100110011100",
            669 => "001100110011100",
            670 => "001100110011100",
            671 => "001100110011100",
            672 => "001101000011000",
            673 => "001101000011000",
            674 => "001101000011000",
            675 => "001101000011000",
            676 => "001101000011000",
            677 => "001101000011000",
            678 => "001101000011000",
            679 => "001101000011000",
            680 => "001101010011111",
            681 => "001101010011111",
            682 => "001101010011111",
            683 => "001101010011111",
            684 => "001101010011111",
            685 => "001101010011111",
            686 => "001101010011111",
            687 => "001101010011111",
            688 => "001101100010001",
            689 => "001101100010001",
            690 => "001101100010001",
            691 => "001101100010001",
            692 => "001101100010001",
            693 => "001101100010001",
            694 => "001101100010001",
            695 => "001101100010001",
            696 => "001101110010110",
            697 => "001101110010110",
            698 => "001101110010110",
            699 => "001101110010110",
            700 => "001101110010110",
            701 => "001101110010110",
            702 => "001101110010110",
            703 => "001101110010110",
            704 => "001110000011001",
            705 => "001110000011001",
            706 => "001110000011001",
            707 => "001110000011001",
            708 => "001110000011001",
            709 => "001110000011001",
            710 => "001110000011001",
            711 => "001110000011001",
            712 => "001110010011110",
            713 => "001110010011110",
            714 => "001110010011110",
            715 => "001110010011110",
            716 => "001110010011110",
            717 => "001110010011110",
            718 => "001110010011110",
            719 => "001110010011110",
            720 => "001110100010000",
            721 => "001110100010000",
            722 => "001110100010000",
            723 => "001110100010000",
            724 => "001110100010000",
            725 => "001110100010000",
            726 => "001110100010000",
            727 => "001110100010000",
            728 => "001110110010111",
            729 => "001110110010111",
            730 => "001110110010111",
            731 => "001110110010111",
            732 => "001110110010111",
            733 => "001110110010111",
            734 => "001110110010111",
            735 => "001110110010111",
            736 => "001111000010011",
            737 => "001111000010011",
            738 => "001111000010011",
            739 => "001111000010011",
            740 => "001111000010011",
            741 => "001111000010011",
            742 => "001111000010011",
            743 => "001111000010011",
            744 => "001111010010100",
            745 => "001111010010100",
            746 => "001111010010100",
            747 => "001111010010100",
            748 => "001111010010100",
            749 => "001111010010100",
            750 => "001111010010100",
            751 => "001111010010100",
            752 => "001111100011010",
            753 => "001111100011010",
            754 => "001111100011010",
            755 => "001111100011010",
            756 => "001111100011010",
            757 => "001111100011010",
            758 => "001111100011010",
            759 => "001111100011010",
            760 => "001111110011101",
            761 => "001111110011101",
            762 => "001111110011101",
            763 => "001111110011101",
            764 => "001111110011101",
            765 => "001111110011101",
            766 => "001111110011101",
            767 => "001111110011101",
            768 => "010000000011101",
            769 => "010000000011101",
            770 => "010000000011101",
            771 => "010000000011101",
            772 => "010000000011101",
            773 => "010000000011101",
            774 => "010000000011101",
            775 => "010000000011101",
            776 => "010000010011010",
            777 => "010000010011010",
            778 => "010000010011010",
            779 => "010000010011010",
            780 => "010000010011010",
            781 => "010000010011010",
            782 => "010000010011010",
            783 => "010000010011010",
            784 => "010000100010100",
            785 => "010000100010100",
            786 => "010000100010100",
            787 => "010000100010100",
            788 => "010000100010100",
            789 => "010000100010100",
            790 => "010000100010100",
            791 => "010000100010100",
            792 => "010000110010011",
            793 => "010000110010011",
            794 => "010000110010011",
            795 => "010000110010011",
            796 => "010000110010011",
            797 => "010000110010011",
            798 => "010000110010011",
            799 => "010000110010011",
            800 => "010001000010111",
            801 => "010001000010111",
            802 => "010001000010111",
            803 => "010001000010111",
            804 => "010001000010111",
            805 => "010001000010111",
            806 => "010001000010111",
            807 => "010001000010111",
            808 => "010001010010000",
            809 => "010001010010000",
            810 => "010001010010000",
            811 => "010001010010000",
            812 => "010001010010000",
            813 => "010001010010000",
            814 => "010001010010000",
            815 => "010001010010000",
            816 => "010001100011110",
            817 => "010001100011110",
            818 => "010001100011110",
            819 => "010001100011110",
            820 => "010001100011110",
            821 => "010001100011110",
            822 => "010001100011110",
            823 => "010001100011110",
            824 => "010001110011001",
            825 => "010001110011001",
            826 => "010001110011001",
            827 => "010001110011001",
            828 => "010001110011001",
            829 => "010001110011001",
            830 => "010001110011001",
            831 => "010001110011001",
            832 => "010010000010110",
            833 => "010010000010110",
            834 => "010010000010110",
            835 => "010010000010110",
            836 => "010010000010110",
            837 => "010010000010110",
            838 => "010010000010110",
            839 => "010010000010110",
            840 => "010010010010001",
            841 => "010010010010001",
            842 => "010010010010001",
            843 => "010010010010001",
            844 => "010010010010001",
            845 => "010010010010001",
            846 => "010010010010001",
            847 => "010010010010001",
            848 => "010010100011111",
            849 => "010010100011111",
            850 => "010010100011111",
            851 => "010010100011111",
            852 => "010010100011111",
            853 => "010010100011111",
            854 => "010010100011111",
            855 => "010010100011111",
            856 => "010010110011000",
            857 => "010010110011000",
            858 => "010010110011000",
            859 => "010010110011000",
            860 => "010010110011000",
            861 => "010010110011000",
            862 => "010010110011000",
            863 => "010010110011000",
            864 => "010011000011100",
            865 => "010011000011100",
            866 => "010011000011100",
            867 => "010011000011100",
            868 => "010011000011100",
            869 => "010011000011100",
            870 => "010011000011100",
            871 => "010011000011100",
            872 => "010011010011011",
            873 => "010011010011011",
            874 => "010011010011011",
            875 => "010011010011011",
            876 => "010011010011011",
            877 => "010011010011011",
            878 => "010011010011011",
            879 => "010011010011011",
            880 => "010011100010101",
            881 => "010011100010101",
            882 => "010011100010101",
            883 => "010011100010101",
            884 => "010011100010101",
            885 => "010011100010101",
            886 => "010011100010101",
            887 => "010011100010101",
            888 => "010011110010010",
            889 => "010011110010010",
            890 => "010011110010010",
            891 => "010011110010010",
            892 => "010011110010010",
            893 => "010011110010010",
            894 => "010011110010010",
            895 => "010011110010010",
            896 => "010100000010001",
            897 => "010100000010001",
            898 => "010100000010001",
            899 => "010100000010001",
            900 => "010100000010001",
            901 => "010100000010001",
            902 => "010100000010001",
            903 => "010100000010001",
            904 => "010100010010110",
            905 => "010100010010110",
            906 => "010100010010110",
            907 => "010100010010110",
            908 => "010100010010110",
            909 => "010100010010110",
            910 => "010100010010110",
            911 => "010100010010110",
            912 => "010100100011000",
            913 => "010100100011000",
            914 => "010100100011000",
            915 => "010100100011000",
            916 => "010100100011000",
            917 => "010100100011000",
            918 => "010100100011000",
            919 => "010100100011000",
            920 => "010100110011111",
            921 => "010100110011111",
            922 => "010100110011111",
            923 => "010100110011111",
            924 => "010100110011111",
            925 => "010100110011111",
            926 => "010100110011111",
            927 => "010100110011111",
            928 => "010101000011011",
            929 => "010101000011011",
            930 => "010101000011011",
            931 => "010101000011011",
            932 => "010101000011011",
            933 => "010101000011011",
            934 => "010101000011011",
            935 => "010101000011011",
            936 => "010101010011100",
            937 => "010101010011100",
            938 => "010101010011100",
            939 => "010101010011100",
            940 => "010101010011100",
            941 => "010101010011100",
            942 => "010101010011100",
            943 => "010101010011100",
            944 => "010101100010010",
            945 => "010101100010010",
            946 => "010101100010010",
            947 => "010101100010010",
            948 => "010101100010010",
            949 => "010101100010010",
            950 => "010101100010010",
            951 => "010101100010010",
            952 => "010101110010101",
            953 => "010101110010101",
            954 => "010101110010101",
            955 => "010101110010101",
            956 => "010101110010101",
            957 => "010101110010101",
            958 => "010101110010101",
            959 => "010101110010101",
            960 => "010110000011010",
            961 => "010110000011010",
            962 => "010110000011010",
            963 => "010110000011010",
            964 => "010110000011010",
            965 => "010110000011010",
            966 => "010110000011010",
            967 => "010110000011010",
            968 => "010110010011101",
            969 => "010110010011101",
            970 => "010110010011101",
            971 => "010110010011101",
            972 => "010110010011101",
            973 => "010110010011101",
            974 => "010110010011101",
            975 => "010110010011101",
            976 => "010110100010011",
            977 => "010110100010011",
            978 => "010110100010011",
            979 => "010110100010011",
            980 => "010110100010011",
            981 => "010110100010011",
            982 => "010110100010011",
            983 => "010110100010011",
            984 => "010110110010100",
            985 => "010110110010100",
            986 => "010110110010100",
            987 => "010110110010100",
            988 => "010110110010100",
            989 => "010110110010100",
            990 => "010110110010100",
            991 => "010110110010100",
            992 => "010111000010000",
            993 => "010111000010000",
            994 => "010111000010000",
            995 => "010111000010000",
            996 => "010111000010000",
            997 => "010111000010000",
            998 => "010111000010000",
            999 => "010111000010000",
            1000 => "010111010010111",
            1001 => "010111010010111",
            1002 => "010111010010111",
            1003 => "010111010010111",
            1004 => "010111010010111",
            1005 => "010111010010111",
            1006 => "010111010010111",
            1007 => "010111010010111",
            1008 => "010111100011001",
            1009 => "010111100011001",
            1010 => "010111100011001",
            1011 => "010111100011001",
            1012 => "010111100011001",
            1013 => "010111100011001",
            1014 => "010111100011001",
            1015 => "010111100011001",
            1016 => "010111110011110",
            1017 => "010111110011110",
            1018 => "010111110011110",
            1019 => "010111110011110",
            1020 => "010111110011110",
            1021 => "010111110011110",
            1022 => "010111110011110",
            1023 => "010111110011110",
            1024 => "011000000010000",
            1025 => "011000000010000",
            1026 => "011000000010000",
            1027 => "011000000010000",
            1028 => "011000000010000",
            1029 => "011000000010000",
            1030 => "011000000010000",
            1031 => "011000000010000",
            1032 => "011000010010111",
            1033 => "011000010010111",
            1034 => "011000010010111",
            1035 => "011000010010111",
            1036 => "011000010010111",
            1037 => "011000010010111",
            1038 => "011000010010111",
            1039 => "011000010010111",
            1040 => "011000100011001",
            1041 => "011000100011001",
            1042 => "011000100011001",
            1043 => "011000100011001",
            1044 => "011000100011001",
            1045 => "011000100011001",
            1046 => "011000100011001",
            1047 => "011000100011001",
            1048 => "011000110011110",
            1049 => "011000110011110",
            1050 => "011000110011110",
            1051 => "011000110011110",
            1052 => "011000110011110",
            1053 => "011000110011110",
            1054 => "011000110011110",
            1055 => "011000110011110",
            1056 => "011001000011010",
            1057 => "011001000011010",
            1058 => "011001000011010",
            1059 => "011001000011010",
            1060 => "011001000011010",
            1061 => "011001000011010",
            1062 => "011001000011010",
            1063 => "011001000011010",
            1064 => "011001010011101",
            1065 => "011001010011101",
            1066 => "011001010011101",
            1067 => "011001010011101",
            1068 => "011001010011101",
            1069 => "011001010011101",
            1070 => "011001010011101",
            1071 => "011001010011101",
            1072 => "011001100010011",
            1073 => "011001100010011",
            1074 => "011001100010011",
            1075 => "011001100010011",
            1076 => "011001100010011",
            1077 => "011001100010011",
            1078 => "011001100010011",
            1079 => "011001100010011",
            1080 => "011001110010100",
            1081 => "011001110010100",
            1082 => "011001110010100",
            1083 => "011001110010100",
            1084 => "011001110010100",
            1085 => "011001110010100",
            1086 => "011001110010100",
            1087 => "011001110010100",
            1088 => "011010000011011",
            1089 => "011010000011011",
            1090 => "011010000011011",
            1091 => "011010000011011",
            1092 => "011010000011011",
            1093 => "011010000011011",
            1094 => "011010000011011",
            1095 => "011010000011011",
            1096 => "011010010011100",
            1097 => "011010010011100",
            1098 => "011010010011100",
            1099 => "011010010011100",
            1100 => "011010010011100",
            1101 => "011010010011100",
            1102 => "011010010011100",
            1103 => "011010010011100",
            1104 => "011010100010010",
            1105 => "011010100010010",
            1106 => "011010100010010",
            1107 => "011010100010010",
            1108 => "011010100010010",
            1109 => "011010100010010",
            1110 => "011010100010010",
            1111 => "011010100010010",
            1112 => "011010110010101",
            1113 => "011010110010101",
            1114 => "011010110010101",
            1115 => "011010110010101",
            1116 => "011010110010101",
            1117 => "011010110010101",
            1118 => "011010110010101",
            1119 => "011010110010101",
            1120 => "011011000010001",
            1121 => "011011000010001",
            1122 => "011011000010001",
            1123 => "011011000010001",
            1124 => "011011000010001",
            1125 => "011011000010001",
            1126 => "011011000010001",
            1127 => "011011000010001",
            1128 => "011011010010110",
            1129 => "011011010010110",
            1130 => "011011010010110",
            1131 => "011011010010110",
            1132 => "011011010010110",
            1133 => "011011010010110",
            1134 => "011011010010110",
            1135 => "011011010010110",
            1136 => "011011100011000",
            1137 => "011011100011000",
            1138 => "011011100011000",
            1139 => "011011100011000",
            1140 => "011011100011000",
            1141 => "011011100011000",
            1142 => "011011100011000",
            1143 => "011011100011000",
            1144 => "011011110011111",
            1145 => "011011110011111",
            1146 => "011011110011111",
            1147 => "011011110011111",
            1148 => "011011110011111",
            1149 => "011011110011111",
            1150 => "011011110011111",
            1151 => "011011110011111",
            1152 => "011100000011100",
            1153 => "011100000011100",
            1154 => "011100000011100",
            1155 => "011100000011100",
            1156 => "011100000011100",
            1157 => "011100000011100",
            1158 => "011100000011100",
            1159 => "011100000011100",
            1160 => "011100010011011",
            1161 => "011100010011011",
            1162 => "011100010011011",
            1163 => "011100010011011",
            1164 => "011100010011011",
            1165 => "011100010011011",
            1166 => "011100010011011",
            1167 => "011100010011011",
            1168 => "011100100010101",
            1169 => "011100100010101",
            1170 => "011100100010101",
            1171 => "011100100010101",
            1172 => "011100100010101",
            1173 => "011100100010101",
            1174 => "011100100010101",
            1175 => "011100100010101",
            1176 => "011100110010010",
            1177 => "011100110010010",
            1178 => "011100110010010",
            1179 => "011100110010010",
            1180 => "011100110010010",
            1181 => "011100110010010",
            1182 => "011100110010010",
            1183 => "011100110010010",
            1184 => "011101000010110",
            1185 => "011101000010110",
            1186 => "011101000010110",
            1187 => "011101000010110",
            1188 => "011101000010110",
            1189 => "011101000010110",
            1190 => "011101000010110",
            1191 => "011101000010110",
            1192 => "011101010010001",
            1193 => "011101010010001",
            1194 => "011101010010001",
            1195 => "011101010010001",
            1196 => "011101010010001",
            1197 => "011101010010001",
            1198 => "011101010010001",
            1199 => "011101010010001",
            1200 => "011101100011111",
            1201 => "011101100011111",
            1202 => "011101100011111",
            1203 => "011101100011111",
            1204 => "011101100011111",
            1205 => "011101100011111",
            1206 => "011101100011111",
            1207 => "011101100011111",
            1208 => "011101110011000",
            1209 => "011101110011000",
            1210 => "011101110011000",
            1211 => "011101110011000",
            1212 => "011101110011000",
            1213 => "011101110011000",
            1214 => "011101110011000",
            1215 => "011101110011000",
            1216 => "011110000010111",
            1217 => "011110000010111",
            1218 => "011110000010111",
            1219 => "011110000010111",
            1220 => "011110000010111",
            1221 => "011110000010111",
            1222 => "011110000010111",
            1223 => "011110000010111",
            1224 => "011110010010000",
            1225 => "011110010010000",
            1226 => "011110010010000",
            1227 => "011110010010000",
            1228 => "011110010010000",
            1229 => "011110010010000",
            1230 => "011110010010000",
            1231 => "011110010010000",
            1232 => "011110100011110",
            1233 => "011110100011110",
            1234 => "011110100011110",
            1235 => "011110100011110",
            1236 => "011110100011110",
            1237 => "011110100011110",
            1238 => "011110100011110",
            1239 => "011110100011110",
            1240 => "011110110011001",
            1241 => "011110110011001",
            1242 => "011110110011001",
            1243 => "011110110011001",
            1244 => "011110110011001",
            1245 => "011110110011001",
            1246 => "011110110011001",
            1247 => "011110110011001",
            1248 => "011111000011101",
            1249 => "011111000011101",
            1250 => "011111000011101",
            1251 => "011111000011101",
            1252 => "011111000011101",
            1253 => "011111000011101",
            1254 => "011111000011101",
            1255 => "011111000011101",
            1256 => "011111010011010",
            1257 => "011111010011010",
            1258 => "011111010011010",
            1259 => "011111010011010",
            1260 => "011111010011010",
            1261 => "011111010011010",
            1262 => "011111010011010",
            1263 => "011111010011010",
            1264 => "011111100010100",
            1265 => "011111100010100",
            1266 => "011111100010100",
            1267 => "011111100010100",
            1268 => "011111100010100",
            1269 => "011111100010100",
            1270 => "011111100010100",
            1271 => "011111100010100",
            1272 => "011111110010011",
            1273 => "011111110010011",
            1274 => "011111110010011",
            1275 => "011111110010011",
            1276 => "011111110010011",
            1277 => "011111110010011",
            1278 => "011111110010011",
            1279 => "011111110010011",
            1280 => "100000000011100",
            1281 => "100000000011100",
            1282 => "100000000011100",
            1283 => "100000000011100",
            1284 => "100000000011100",
            1285 => "100000000011100",
            1286 => "100000000011100",
            1287 => "100000000011100",
            1288 => "100000010011011",
            1289 => "100000010011011",
            1290 => "100000010011011",
            1291 => "100000010011011",
            1292 => "100000010011011",
            1293 => "100000010011011",
            1294 => "100000010011011",
            1295 => "100000010011011",
            1296 => "100000100010101",
            1297 => "100000100010101",
            1298 => "100000100010101",
            1299 => "100000100010101",
            1300 => "100000100010101",
            1301 => "100000100010101",
            1302 => "100000100010101",
            1303 => "100000100010101",
            1304 => "100000110010010",
            1305 => "100000110010010",
            1306 => "100000110010010",
            1307 => "100000110010010",
            1308 => "100000110010010",
            1309 => "100000110010010",
            1310 => "100000110010010",
            1311 => "100000110010010",
            1312 => "100001000010110",
            1313 => "100001000010110",
            1314 => "100001000010110",
            1315 => "100001000010110",
            1316 => "100001000010110",
            1317 => "100001000010110",
            1318 => "100001000010110",
            1319 => "100001000010110",
            1320 => "100001010010001",
            1321 => "100001010010001",
            1322 => "100001010010001",
            1323 => "100001010010001",
            1324 => "100001010010001",
            1325 => "100001010010001",
            1326 => "100001010010001",
            1327 => "100001010010001",
            1328 => "100001100011111",
            1329 => "100001100011111",
            1330 => "100001100011111",
            1331 => "100001100011111",
            1332 => "100001100011111",
            1333 => "100001100011111",
            1334 => "100001100011111",
            1335 => "100001100011111",
            1336 => "100001110011000",
            1337 => "100001110011000",
            1338 => "100001110011000",
            1339 => "100001110011000",
            1340 => "100001110011000",
            1341 => "100001110011000",
            1342 => "100001110011000",
            1343 => "100001110011000",
            1344 => "100010000010111",
            1345 => "100010000010111",
            1346 => "100010000010111",
            1347 => "100010000010111",
            1348 => "100010000010111",
            1349 => "100010000010111",
            1350 => "100010000010111",
            1351 => "100010000010111",
            1352 => "100010010010000",
            1353 => "100010010010000",
            1354 => "100010010010000",
            1355 => "100010010010000",
            1356 => "100010010010000",
            1357 => "100010010010000",
            1358 => "100010010010000",
            1359 => "100010010010000",
            1360 => "100010100011110",
            1361 => "100010100011110",
            1362 => "100010100011110",
            1363 => "100010100011110",
            1364 => "100010100011110",
            1365 => "100010100011110",
            1366 => "100010100011110",
            1367 => "100010100011110",
            1368 => "100010110011001",
            1369 => "100010110011001",
            1370 => "100010110011001",
            1371 => "100010110011001",
            1372 => "100010110011001",
            1373 => "100010110011001",
            1374 => "100010110011001",
            1375 => "100010110011001",
            1376 => "100011000011101",
            1377 => "100011000011101",
            1378 => "100011000011101",
            1379 => "100011000011101",
            1380 => "100011000011101",
            1381 => "100011000011101",
            1382 => "100011000011101",
            1383 => "100011000011101",
            1384 => "100011010011010",
            1385 => "100011010011010",
            1386 => "100011010011010",
            1387 => "100011010011010",
            1388 => "100011010011010",
            1389 => "100011010011010",
            1390 => "100011010011010",
            1391 => "100011010011010",
            1392 => "100011100010100",
            1393 => "100011100010100",
            1394 => "100011100010100",
            1395 => "100011100010100",
            1396 => "100011100010100",
            1397 => "100011100010100",
            1398 => "100011100010100",
            1399 => "100011100010100",
            1400 => "100011110010011",
            1401 => "100011110010011",
            1402 => "100011110010011",
            1403 => "100011110010011",
            1404 => "100011110010011",
            1405 => "100011110010011",
            1406 => "100011110010011",
            1407 => "100011110010011",
            1408 => "100100000010000",
            1409 => "100100000010000",
            1410 => "100100000010000",
            1411 => "100100000010000",
            1412 => "100100000010000",
            1413 => "100100000010000",
            1414 => "100100000010000",
            1415 => "100100000010000",
            1416 => "100100010010111",
            1417 => "100100010010111",
            1418 => "100100010010111",
            1419 => "100100010010111",
            1420 => "100100010010111",
            1421 => "100100010010111",
            1422 => "100100010010111",
            1423 => "100100010010111",
            1424 => "100100100011001",
            1425 => "100100100011001",
            1426 => "100100100011001",
            1427 => "100100100011001",
            1428 => "100100100011001",
            1429 => "100100100011001",
            1430 => "100100100011001",
            1431 => "100100100011001",
            1432 => "100100110011110",
            1433 => "100100110011110",
            1434 => "100100110011110",
            1435 => "100100110011110",
            1436 => "100100110011110",
            1437 => "100100110011110",
            1438 => "100100110011110",
            1439 => "100100110011110",
            1440 => "100101000011010",
            1441 => "100101000011010",
            1442 => "100101000011010",
            1443 => "100101000011010",
            1444 => "100101000011010",
            1445 => "100101000011010",
            1446 => "100101000011010",
            1447 => "100101000011010",
            1448 => "100101010011101",
            1449 => "100101010011101",
            1450 => "100101010011101",
            1451 => "100101010011101",
            1452 => "100101010011101",
            1453 => "100101010011101",
            1454 => "100101010011101",
            1455 => "100101010011101",
            1456 => "100101100010011",
            1457 => "100101100010011",
            1458 => "100101100010011",
            1459 => "100101100010011",
            1460 => "100101100010011",
            1461 => "100101100010011",
            1462 => "100101100010011",
            1463 => "100101100010011",
            1464 => "100101110010100",
            1465 => "100101110010100",
            1466 => "100101110010100",
            1467 => "100101110010100",
            1468 => "100101110010100",
            1469 => "100101110010100",
            1470 => "100101110010100",
            1471 => "100101110010100",
            1472 => "100110000011011",
            1473 => "100110000011011",
            1474 => "100110000011011",
            1475 => "100110000011011",
            1476 => "100110000011011",
            1477 => "100110000011011",
            1478 => "100110000011011",
            1479 => "100110000011011",
            1480 => "100110010011100",
            1481 => "100110010011100",
            1482 => "100110010011100",
            1483 => "100110010011100",
            1484 => "100110010011100",
            1485 => "100110010011100",
            1486 => "100110010011100",
            1487 => "100110010011100",
            1488 => "100110100010010",
            1489 => "100110100010010",
            1490 => "100110100010010",
            1491 => "100110100010010",
            1492 => "100110100010010",
            1493 => "100110100010010",
            1494 => "100110100010010",
            1495 => "100110100010010",
            1496 => "100110110010101",
            1497 => "100110110010101",
            1498 => "100110110010101",
            1499 => "100110110010101",
            1500 => "100110110010101",
            1501 => "100110110010101",
            1502 => "100110110010101",
            1503 => "100110110010101",
            1504 => "100111000010001",
            1505 => "100111000010001",
            1506 => "100111000010001",
            1507 => "100111000010001",
            1508 => "100111000010001",
            1509 => "100111000010001",
            1510 => "100111000010001",
            1511 => "100111000010001",
            1512 => "100111010010110",
            1513 => "100111010010110",
            1514 => "100111010010110",
            1515 => "100111010010110",
            1516 => "100111010010110",
            1517 => "100111010010110",
            1518 => "100111010010110",
            1519 => "100111010010110",
            1520 => "100111100011000",
            1521 => "100111100011000",
            1522 => "100111100011000",
            1523 => "100111100011000",
            1524 => "100111100011000",
            1525 => "100111100011000",
            1526 => "100111100011000",
            1527 => "100111100011000",
            1528 => "100111110011111",
            1529 => "100111110011111",
            1530 => "100111110011111",
            1531 => "100111110011111",
            1532 => "100111110011111",
            1533 => "100111110011111",
            1534 => "100111110011111",
            1535 => "100111110011111",
            1536 => "101000000010001",
            1537 => "101000000010001",
            1538 => "101000000010001",
            1539 => "101000000010001",
            1540 => "101000000010001",
            1541 => "101000000010001",
            1542 => "101000000010001",
            1543 => "101000000010001",
            1544 => "101000010010110",
            1545 => "101000010010110",
            1546 => "101000010010110",
            1547 => "101000010010110",
            1548 => "101000010010110",
            1549 => "101000010010110",
            1550 => "101000010010110",
            1551 => "101000010010110",
            1552 => "101000100011000",
            1553 => "101000100011000",
            1554 => "101000100011000",
            1555 => "101000100011000",
            1556 => "101000100011000",
            1557 => "101000100011000",
            1558 => "101000100011000",
            1559 => "101000100011000",
            1560 => "101000110011111",
            1561 => "101000110011111",
            1562 => "101000110011111",
            1563 => "101000110011111",
            1564 => "101000110011111",
            1565 => "101000110011111",
            1566 => "101000110011111",
            1567 => "101000110011111",
            1568 => "101001000011011",
            1569 => "101001000011011",
            1570 => "101001000011011",
            1571 => "101001000011011",
            1572 => "101001000011011",
            1573 => "101001000011011",
            1574 => "101001000011011",
            1575 => "101001000011011",
            1576 => "101001010011100",
            1577 => "101001010011100",
            1578 => "101001010011100",
            1579 => "101001010011100",
            1580 => "101001010011100",
            1581 => "101001010011100",
            1582 => "101001010011100",
            1583 => "101001010011100",
            1584 => "101001100010010",
            1585 => "101001100010010",
            1586 => "101001100010010",
            1587 => "101001100010010",
            1588 => "101001100010010",
            1589 => "101001100010010",
            1590 => "101001100010010",
            1591 => "101001100010010",
            1592 => "101001110010101",
            1593 => "101001110010101",
            1594 => "101001110010101",
            1595 => "101001110010101",
            1596 => "101001110010101",
            1597 => "101001110010101",
            1598 => "101001110010101",
            1599 => "101001110010101",
            1600 => "101010000011010",
            1601 => "101010000011010",
            1602 => "101010000011010",
            1603 => "101010000011010",
            1604 => "101010000011010",
            1605 => "101010000011010",
            1606 => "101010000011010",
            1607 => "101010000011010",
            1608 => "101010010011101",
            1609 => "101010010011101",
            1610 => "101010010011101",
            1611 => "101010010011101",
            1612 => "101010010011101",
            1613 => "101010010011101",
            1614 => "101010010011101",
            1615 => "101010010011101",
            1616 => "101010100010011",
            1617 => "101010100010011",
            1618 => "101010100010011",
            1619 => "101010100010011",
            1620 => "101010100010011",
            1621 => "101010100010011",
            1622 => "101010100010011",
            1623 => "101010100010011",
            1624 => "101010110010100",
            1625 => "101010110010100",
            1626 => "101010110010100",
            1627 => "101010110010100",
            1628 => "101010110010100",
            1629 => "101010110010100",
            1630 => "101010110010100",
            1631 => "101010110010100",
            1632 => "101011000010000",
            1633 => "101011000010000",
            1634 => "101011000010000",
            1635 => "101011000010000",
            1636 => "101011000010000",
            1637 => "101011000010000",
            1638 => "101011000010000",
            1639 => "101011000010000",
            1640 => "101011010010111",
            1641 => "101011010010111",
            1642 => "101011010010111",
            1643 => "101011010010111",
            1644 => "101011010010111",
            1645 => "101011010010111",
            1646 => "101011010010111",
            1647 => "101011010010111",
            1648 => "101011100011001",
            1649 => "101011100011001",
            1650 => "101011100011001",
            1651 => "101011100011001",
            1652 => "101011100011001",
            1653 => "101011100011001",
            1654 => "101011100011001",
            1655 => "101011100011001",
            1656 => "101011110011110",
            1657 => "101011110011110",
            1658 => "101011110011110",
            1659 => "101011110011110",
            1660 => "101011110011110",
            1661 => "101011110011110",
            1662 => "101011110011110",
            1663 => "101011110011110",
            1664 => "101100000011101",
            1665 => "101100000011101",
            1666 => "101100000011101",
            1667 => "101100000011101",
            1668 => "101100000011101",
            1669 => "101100000011101",
            1670 => "101100000011101",
            1671 => "101100000011101",
            1672 => "101100010011010",
            1673 => "101100010011010",
            1674 => "101100010011010",
            1675 => "101100010011010",
            1676 => "101100010011010",
            1677 => "101100010011010",
            1678 => "101100010011010",
            1679 => "101100010011010",
            1680 => "101100100010100",
            1681 => "101100100010100",
            1682 => "101100100010100",
            1683 => "101100100010100",
            1684 => "101100100010100",
            1685 => "101100100010100",
            1686 => "101100100010100",
            1687 => "101100100010100",
            1688 => "101100110010011",
            1689 => "101100110010011",
            1690 => "101100110010011",
            1691 => "101100110010011",
            1692 => "101100110010011",
            1693 => "101100110010011",
            1694 => "101100110010011",
            1695 => "101100110010011",
            1696 => "101101000010111",
            1697 => "101101000010111",
            1698 => "101101000010111",
            1699 => "101101000010111",
            1700 => "101101000010111",
            1701 => "101101000010111",
            1702 => "101101000010111",
            1703 => "101101000010111",
            1704 => "101101010010000",
            1705 => "101101010010000",
            1706 => "101101010010000",
            1707 => "101101010010000",
            1708 => "101101010010000",
            1709 => "101101010010000",
            1710 => "101101010010000",
            1711 => "101101010010000",
            1712 => "101101100011110",
            1713 => "101101100011110",
            1714 => "101101100011110",
            1715 => "101101100011110",
            1716 => "101101100011110",
            1717 => "101101100011110",
            1718 => "101101100011110",
            1719 => "101101100011110",
            1720 => "101101110011001",
            1721 => "101101110011001",
            1722 => "101101110011001",
            1723 => "101101110011001",
            1724 => "101101110011001",
            1725 => "101101110011001",
            1726 => "101101110011001",
            1727 => "101101110011001",
            1728 => "101110000010110",
            1729 => "101110000010110",
            1730 => "101110000010110",
            1731 => "101110000010110",
            1732 => "101110000010110",
            1733 => "101110000010110",
            1734 => "101110000010110",
            1735 => "101110000010110",
            1736 => "101110010010001",
            1737 => "101110010010001",
            1738 => "101110010010001",
            1739 => "101110010010001",
            1740 => "101110010010001",
            1741 => "101110010010001",
            1742 => "101110010010001",
            1743 => "101110010010001",
            1744 => "101110100011111",
            1745 => "101110100011111",
            1746 => "101110100011111",
            1747 => "101110100011111",
            1748 => "101110100011111",
            1749 => "101110100011111",
            1750 => "101110100011111",
            1751 => "101110100011111",
            1752 => "101110110011000",
            1753 => "101110110011000",
            1754 => "101110110011000",
            1755 => "101110110011000",
            1756 => "101110110011000",
            1757 => "101110110011000",
            1758 => "101110110011000",
            1759 => "101110110011000",
            1760 => "101111000011100",
            1761 => "101111000011100",
            1762 => "101111000011100",
            1763 => "101111000011100",
            1764 => "101111000011100",
            1765 => "101111000011100",
            1766 => "101111000011100",
            1767 => "101111000011100",
            1768 => "101111010011011",
            1769 => "101111010011011",
            1770 => "101111010011011",
            1771 => "101111010011011",
            1772 => "101111010011011",
            1773 => "101111010011011",
            1774 => "101111010011011",
            1775 => "101111010011011",
            1776 => "101111100010101",
            1777 => "101111100010101",
            1778 => "101111100010101",
            1779 => "101111100010101",
            1780 => "101111100010101",
            1781 => "101111100010101",
            1782 => "101111100010101",
            1783 => "101111100010101",
            1784 => "101111110010010",
            1785 => "101111110010010",
            1786 => "101111110010010",
            1787 => "101111110010010",
            1788 => "101111110010010",
            1789 => "101111110010010",
            1790 => "101111110010010",
            1791 => "101111110010010",
            1792 => "110000000010010",
            1793 => "110000000010010",
            1794 => "110000000010010",
            1795 => "110000000010010",
            1796 => "110000000010010",
            1797 => "110000000010010",
            1798 => "110000000010010",
            1799 => "110000000010010",
            1800 => "110000010010101",
            1801 => "110000010010101",
            1802 => "110000010010101",
            1803 => "110000010010101",
            1804 => "110000010010101",
            1805 => "110000010010101",
            1806 => "110000010010101",
            1807 => "110000010010101",
            1808 => "110000100011011",
            1809 => "110000100011011",
            1810 => "110000100011011",
            1811 => "110000100011011",
            1812 => "110000100011011",
            1813 => "110000100011011",
            1814 => "110000100011011",
            1815 => "110000100011011",
            1816 => "110000110011100",
            1817 => "110000110011100",
            1818 => "110000110011100",
            1819 => "110000110011100",
            1820 => "110000110011100",
            1821 => "110000110011100",
            1822 => "110000110011100",
            1823 => "110000110011100",
            1824 => "110001000011000",
            1825 => "110001000011000",
            1826 => "110001000011000",
            1827 => "110001000011000",
            1828 => "110001000011000",
            1829 => "110001000011000",
            1830 => "110001000011000",
            1831 => "110001000011000",
            1832 => "110001010011111",
            1833 => "110001010011111",
            1834 => "110001010011111",
            1835 => "110001010011111",
            1836 => "110001010011111",
            1837 => "110001010011111",
            1838 => "110001010011111",
            1839 => "110001010011111",
            1840 => "110001100010001",
            1841 => "110001100010001",
            1842 => "110001100010001",
            1843 => "110001100010001",
            1844 => "110001100010001",
            1845 => "110001100010001",
            1846 => "110001100010001",
            1847 => "110001100010001",
            1848 => "110001110010110",
            1849 => "110001110010110",
            1850 => "110001110010110",
            1851 => "110001110010110",
            1852 => "110001110010110",
            1853 => "110001110010110",
            1854 => "110001110010110",
            1855 => "110001110010110",
            1856 => "110010000011001",
            1857 => "110010000011001",
            1858 => "110010000011001",
            1859 => "110010000011001",
            1860 => "110010000011001",
            1861 => "110010000011001",
            1862 => "110010000011001",
            1863 => "110010000011001",
            1864 => "110010010011110",
            1865 => "110010010011110",
            1866 => "110010010011110",
            1867 => "110010010011110",
            1868 => "110010010011110",
            1869 => "110010010011110",
            1870 => "110010010011110",
            1871 => "110010010011110",
            1872 => "110010100010000",
            1873 => "110010100010000",
            1874 => "110010100010000",
            1875 => "110010100010000",
            1876 => "110010100010000",
            1877 => "110010100010000",
            1878 => "110010100010000",
            1879 => "110010100010000",
            1880 => "110010110010111",
            1881 => "110010110010111",
            1882 => "110010110010111",
            1883 => "110010110010111",
            1884 => "110010110010111",
            1885 => "110010110010111",
            1886 => "110010110010111",
            1887 => "110010110010111",
            1888 => "110011000010011",
            1889 => "110011000010011",
            1890 => "110011000010011",
            1891 => "110011000010011",
            1892 => "110011000010011",
            1893 => "110011000010011",
            1894 => "110011000010011",
            1895 => "110011000010011",
            1896 => "110011010010100",
            1897 => "110011010010100",
            1898 => "110011010010100",
            1899 => "110011010010100",
            1900 => "110011010010100",
            1901 => "110011010010100",
            1902 => "110011010010100",
            1903 => "110011010010100",
            1904 => "110011100011010",
            1905 => "110011100011010",
            1906 => "110011100011010",
            1907 => "110011100011010",
            1908 => "110011100011010",
            1909 => "110011100011010",
            1910 => "110011100011010",
            1911 => "110011100011010",
            1912 => "110011110011101",
            1913 => "110011110011101",
            1914 => "110011110011101",
            1915 => "110011110011101",
            1916 => "110011110011101",
            1917 => "110011110011101",
            1918 => "110011110011101",
            1919 => "110011110011101",
            1920 => "110100000011110",
            1921 => "110100000011110",
            1922 => "110100000011110",
            1923 => "110100000011110",
            1924 => "110100000011110",
            1925 => "110100000011110",
            1926 => "110100000011110",
            1927 => "110100000011110",
            1928 => "110100010011001",
            1929 => "110100010011001",
            1930 => "110100010011001",
            1931 => "110100010011001",
            1932 => "110100010011001",
            1933 => "110100010011001",
            1934 => "110100010011001",
            1935 => "110100010011001",
            1936 => "110100100010111",
            1937 => "110100100010111",
            1938 => "110100100010111",
            1939 => "110100100010111",
            1940 => "110100100010111",
            1941 => "110100100010111",
            1942 => "110100100010111",
            1943 => "110100100010111",
            1944 => "110100110010000",
            1945 => "110100110010000",
            1946 => "110100110010000",
            1947 => "110100110010000",
            1948 => "110100110010000",
            1949 => "110100110010000",
            1950 => "110100110010000",
            1951 => "110100110010000",
            1952 => "110101000010100",
            1953 => "110101000010100",
            1954 => "110101000010100",
            1955 => "110101000010100",
            1956 => "110101000010100",
            1957 => "110101000010100",
            1958 => "110101000010100",
            1959 => "110101000010100",
            1960 => "110101010010011",
            1961 => "110101010010011",
            1962 => "110101010010011",
            1963 => "110101010010011",
            1964 => "110101010010011",
            1965 => "110101010010011",
            1966 => "110101010010011",
            1967 => "110101010010011",
            1968 => "110101100011101",
            1969 => "110101100011101",
            1970 => "110101100011101",
            1971 => "110101100011101",
            1972 => "110101100011101",
            1973 => "110101100011101",
            1974 => "110101100011101",
            1975 => "110101100011101",
            1976 => "110101110011010",
            1977 => "110101110011010",
            1978 => "110101110011010",
            1979 => "110101110011010",
            1980 => "110101110011010",
            1981 => "110101110011010",
            1982 => "110101110011010",
            1983 => "110101110011010",
            1984 => "110110000010101",
            1985 => "110110000010101",
            1986 => "110110000010101",
            1987 => "110110000010101",
            1988 => "110110000010101",
            1989 => "110110000010101",
            1990 => "110110000010101",
            1991 => "110110000010101",
            1992 => "110110010010010",
            1993 => "110110010010010",
            1994 => "110110010010010",
            1995 => "110110010010010",
            1996 => "110110010010010",
            1997 => "110110010010010",
            1998 => "110110010010010",
            1999 => "110110010010010",
            2000 => "110110100011100",
            2001 => "110110100011100",
            2002 => "110110100011100",
            2003 => "110110100011100",
            2004 => "110110100011100",
            2005 => "110110100011100",
            2006 => "110110100011100",
            2007 => "110110100011100",
            2008 => "110110110011011",
            2009 => "110110110011011",
            2010 => "110110110011011",
            2011 => "110110110011011",
            2012 => "110110110011011",
            2013 => "110110110011011",
            2014 => "110110110011011",
            2015 => "110110110011011",
            2016 => "110111000011111",
            2017 => "110111000011111",
            2018 => "110111000011111",
            2019 => "110111000011111",
            2020 => "110111000011111",
            2021 => "110111000011111",
            2022 => "110111000011111",
            2023 => "110111000011111",
            2024 => "110111010011000",
            2025 => "110111010011000",
            2026 => "110111010011000",
            2027 => "110111010011000",
            2028 => "110111010011000",
            2029 => "110111010011000",
            2030 => "110111010011000",
            2031 => "110111010011000",
            2032 => "110111100010110",
            2033 => "110111100010110",
            2034 => "110111100010110",
            2035 => "110111100010110",
            2036 => "110111100010110",
            2037 => "110111100010110",
            2038 => "110111100010110",
            2039 => "110111100010110",
            2040 => "110111110010001",
            2041 => "110111110010001",
            2042 => "110111110010001",
            2043 => "110111110010001",
            2044 => "110111110010001",
            2045 => "110111110010001",
            2046 => "110111110010001",
            2047 => "110111110010001",
            2048 => "111000000011111",
            2049 => "111000000011111",
            2050 => "111000000011111",
            2051 => "111000000011111",
            2052 => "111000000011111",
            2053 => "111000000011111",
            2054 => "111000000011111",
            2055 => "111000000011111",
            2056 => "111000010011000",
            2057 => "111000010011000",
            2058 => "111000010011000",
            2059 => "111000010011000",
            2060 => "111000010011000",
            2061 => "111000010011000",
            2062 => "111000010011000",
            2063 => "111000010011000",
            2064 => "111000100010110",
            2065 => "111000100010110",
            2066 => "111000100010110",
            2067 => "111000100010110",
            2068 => "111000100010110",
            2069 => "111000100010110",
            2070 => "111000100010110",
            2071 => "111000100010110",
            2072 => "111000110010001",
            2073 => "111000110010001",
            2074 => "111000110010001",
            2075 => "111000110010001",
            2076 => "111000110010001",
            2077 => "111000110010001",
            2078 => "111000110010001",
            2079 => "111000110010001",
            2080 => "111001000010101",
            2081 => "111001000010101",
            2082 => "111001000010101",
            2083 => "111001000010101",
            2084 => "111001000010101",
            2085 => "111001000010101",
            2086 => "111001000010101",
            2087 => "111001000010101",
            2088 => "111001010010010",
            2089 => "111001010010010",
            2090 => "111001010010010",
            2091 => "111001010010010",
            2092 => "111001010010010",
            2093 => "111001010010010",
            2094 => "111001010010010",
            2095 => "111001010010010",
            2096 => "111001100011100",
            2097 => "111001100011100",
            2098 => "111001100011100",
            2099 => "111001100011100",
            2100 => "111001100011100",
            2101 => "111001100011100",
            2102 => "111001100011100",
            2103 => "111001100011100",
            2104 => "111001110011011",
            2105 => "111001110011011",
            2106 => "111001110011011",
            2107 => "111001110011011",
            2108 => "111001110011011",
            2109 => "111001110011011",
            2110 => "111001110011011",
            2111 => "111001110011011",
            2112 => "111010000010100",
            2113 => "111010000010100",
            2114 => "111010000010100",
            2115 => "111010000010100",
            2116 => "111010000010100",
            2117 => "111010000010100",
            2118 => "111010000010100",
            2119 => "111010000010100",
            2120 => "111010010010011",
            2121 => "111010010010011",
            2122 => "111010010010011",
            2123 => "111010010010011",
            2124 => "111010010010011",
            2125 => "111010010010011",
            2126 => "111010010010011",
            2127 => "111010010010011",
            2128 => "111010100011101",
            2129 => "111010100011101",
            2130 => "111010100011101",
            2131 => "111010100011101",
            2132 => "111010100011101",
            2133 => "111010100011101",
            2134 => "111010100011101",
            2135 => "111010100011101",
            2136 => "111010110011010",
            2137 => "111010110011010",
            2138 => "111010110011010",
            2139 => "111010110011010",
            2140 => "111010110011010",
            2141 => "111010110011010",
            2142 => "111010110011010",
            2143 => "111010110011010",
            2144 => "111011000011110",
            2145 => "111011000011110",
            2146 => "111011000011110",
            2147 => "111011000011110",
            2148 => "111011000011110",
            2149 => "111011000011110",
            2150 => "111011000011110",
            2151 => "111011000011110",
            2152 => "111011010011001",
            2153 => "111011010011001",
            2154 => "111011010011001",
            2155 => "111011010011001",
            2156 => "111011010011001",
            2157 => "111011010011001",
            2158 => "111011010011001",
            2159 => "111011010011001",
            2160 => "111011100010111",
            2161 => "111011100010111",
            2162 => "111011100010111",
            2163 => "111011100010111",
            2164 => "111011100010111",
            2165 => "111011100010111",
            2166 => "111011100010111",
            2167 => "111011100010111",
            2168 => "111011110010000",
            2169 => "111011110010000",
            2170 => "111011110010000",
            2171 => "111011110010000",
            2172 => "111011110010000",
            2173 => "111011110010000",
            2174 => "111011110010000",
            2175 => "111011110010000",
            2176 => "111100000010011",
            2177 => "111100000010011",
            2178 => "111100000010011",
            2179 => "111100000010011",
            2180 => "111100000010011",
            2181 => "111100000010011",
            2182 => "111100000010011",
            2183 => "111100000010011",
            2184 => "111100010010100",
            2185 => "111100010010100",
            2186 => "111100010010100",
            2187 => "111100010010100",
            2188 => "111100010010100",
            2189 => "111100010010100",
            2190 => "111100010010100",
            2191 => "111100010010100",
            2192 => "111100100011010",
            2193 => "111100100011010",
            2194 => "111100100011010",
            2195 => "111100100011010",
            2196 => "111100100011010",
            2197 => "111100100011010",
            2198 => "111100100011010",
            2199 => "111100100011010",
            2200 => "111100110011101",
            2201 => "111100110011101",
            2202 => "111100110011101",
            2203 => "111100110011101",
            2204 => "111100110011101",
            2205 => "111100110011101",
            2206 => "111100110011101",
            2207 => "111100110011101",
            2208 => "111101000011001",
            2209 => "111101000011001",
            2210 => "111101000011001",
            2211 => "111101000011001",
            2212 => "111101000011001",
            2213 => "111101000011001",
            2214 => "111101000011001",
            2215 => "111101000011001",
            2216 => "111101010011110",
            2217 => "111101010011110",
            2218 => "111101010011110",
            2219 => "111101010011110",
            2220 => "111101010011110",
            2221 => "111101010011110",
            2222 => "111101010011110",
            2223 => "111101010011110",
            2224 => "111101100010000",
            2225 => "111101100010000",
            2226 => "111101100010000",
            2227 => "111101100010000",
            2228 => "111101100010000",
            2229 => "111101100010000",
            2230 => "111101100010000",
            2231 => "111101100010000",
            2232 => "111101110010111",
            2233 => "111101110010111",
            2234 => "111101110010111",
            2235 => "111101110010111",
            2236 => "111101110010111",
            2237 => "111101110010111",
            2238 => "111101110010111",
            2239 => "111101110010111",
            2240 => "111110000011000",
            2241 => "111110000011000",
            2242 => "111110000011000",
            2243 => "111110000011000",
            2244 => "111110000011000",
            2245 => "111110000011000",
            2246 => "111110000011000",
            2247 => "111110000011000",
            2248 => "111110010011111",
            2249 => "111110010011111",
            2250 => "111110010011111",
            2251 => "111110010011111",
            2252 => "111110010011111",
            2253 => "111110010011111",
            2254 => "111110010011111",
            2255 => "111110010011111",
            2256 => "111110100010001",
            2257 => "111110100010001",
            2258 => "111110100010001",
            2259 => "111110100010001",
            2260 => "111110100010001",
            2261 => "111110100010001",
            2262 => "111110100010001",
            2263 => "111110100010001",
            2264 => "111110110010110",
            2265 => "111110110010110",
            2266 => "111110110010110",
            2267 => "111110110010110",
            2268 => "111110110010110",
            2269 => "111110110010110",
            2270 => "111110110010110",
            2271 => "111110110010110",
            2272 => "111111000010010",
            2273 => "111111000010010",
            2274 => "111111000010010",
            2275 => "111111000010010",
            2276 => "111111000010010",
            2277 => "111111000010010",
            2278 => "111111000010010",
            2279 => "111111000010010",
            2280 => "111111010010101",
            2281 => "111111010010101",
            2282 => "111111010010101",
            2283 => "111111010010101",
            2284 => "111111010010101",
            2285 => "111111010010101",
            2286 => "111111010010101",
            2287 => "111111010010101",
            2288 => "111111100011011",
            2289 => "111111100011011",
            2290 => "111111100011011",
            2291 => "111111100011011",
            2292 => "111111100011011",
            2293 => "111111100011011",
            2294 => "111111100011011",
            2295 => "111111100011011",
            2296 => "111111110011100",
            2297 => "111111110011100",
            2298 => "111111110011100",
            2299 => "111111110011100",
            2300 => "111111110011100",
            2301 => "111111110011100",
            2302 => "111111110011100",
            2303 => "111111110011100",
            2304 => "000000000100101",
            2305 => "000000000100101",
            2306 => "000000000100101",
            2307 => "000000000100101",
            2308 => "000000000100101",
            2309 => "000000000100101",
            2310 => "000000000100101",
            2311 => "000000010100010",
            2312 => "000000010100010",
            2313 => "000000010100010",
            2314 => "000000010100010",
            2315 => "000000010100010",
            2316 => "000000010100010",
            2317 => "000000010100010",
            2318 => "000000100101100",
            2319 => "000000100101100",
            2320 => "000000100101100",
            2321 => "000000100101100",
            2322 => "000000100101100",
            2323 => "000000100101100",
            2324 => "000000100101100",
            2325 => "000000110101011",
            2326 => "000000110101011",
            2327 => "000000110101011",
            2328 => "000000110101011",
            2329 => "000000110101011",
            2330 => "000000110101011",
            2331 => "000000110101011",
            2332 => "000001000101111",
            2333 => "000001000101111",
            2334 => "000001000101111",
            2335 => "000001000101111",
            2336 => "000001000101111",
            2337 => "000001000101111",
            2338 => "000001000101111",
            2339 => "000001010101000",
            2340 => "000001010101000",
            2341 => "000001010101000",
            2342 => "000001010101000",
            2343 => "000001010101000",
            2344 => "000001010101000",
            2345 => "000001010101000",
            2346 => "000001100100110",
            2347 => "000001100100110",
            2348 => "000001100100110",
            2349 => "000001100100110",
            2350 => "000001100100110",
            2351 => "000001100100110",
            2352 => "000001100100110",
            2353 => "000001110100001",
            2354 => "000001110100001",
            2355 => "000001110100001",
            2356 => "000001110100001",
            2357 => "000001110100001",
            2358 => "000001110100001",
            2359 => "000001110100001",
            2360 => "000010000101110",
            2361 => "000010000101110",
            2362 => "000010000101110",
            2363 => "000010000101110",
            2364 => "000010000101110",
            2365 => "000010000101110",
            2366 => "000010000101110",
            2367 => "000010010101001",
            2368 => "000010010101001",
            2369 => "000010010101001",
            2370 => "000010010101001",
            2371 => "000010010101001",
            2372 => "000010010101001",
            2373 => "000010010101001",
            2374 => "000010100100111",
            2375 => "000010100100111",
            2376 => "000010100100111",
            2377 => "000010100100111",
            2378 => "000010100100111",
            2379 => "000010100100111",
            2380 => "000010100100111",
            2381 => "000010110100000",
            2382 => "000010110100000",
            2383 => "000010110100000",
            2384 => "000010110100000",
            2385 => "000010110100000",
            2386 => "000010110100000",
            2387 => "000010110100000",
            2388 => "000011000100100",
            2389 => "000011000100100",
            2390 => "000011000100100",
            2391 => "000011000100100",
            2392 => "000011000100100",
            2393 => "000011000100100",
            2394 => "000011000100100",
            2395 => "000011010100011",
            2396 => "000011010100011",
            2397 => "000011010100011",
            2398 => "000011010100011",
            2399 => "000011010100011",
            2400 => "000011010100011",
            2401 => "000011010100011",
            2402 => "000011100101101",
            2403 => "000011100101101",
            2404 => "000011100101101",
            2405 => "000011100101101",
            2406 => "000011100101101",
            2407 => "000011100101101",
            2408 => "000011100101101",
            2409 => "000011110101010",
            2410 => "000011110101010",
            2411 => "000011110101010",
            2412 => "000011110101010",
            2413 => "000011110101010",
            2414 => "000011110101010",
            2415 => "000011110101010",
            2416 => "000100000101001",
            2417 => "000100000101001",
            2418 => "000100000101001",
            2419 => "000100000101001",
            2420 => "000100000101001",
            2421 => "000100000101001",
            2422 => "000100000101001",
            2423 => "000100010101110",
            2424 => "000100010101110",
            2425 => "000100010101110",
            2426 => "000100010101110",
            2427 => "000100010101110",
            2428 => "000100010101110",
            2429 => "000100010101110",
            2430 => "000100100100000",
            2431 => "000100100100000",
            2432 => "000100100100000",
            2433 => "000100100100000",
            2434 => "000100100100000",
            2435 => "000100100100000",
            2436 => "000100100100000",
            2437 => "000100110100111",
            2438 => "000100110100111",
            2439 => "000100110100111",
            2440 => "000100110100111",
            2441 => "000100110100111",
            2442 => "000100110100111",
            2443 => "000100110100111",
            2444 => "000101000100011",
            2445 => "000101000100011",
            2446 => "000101000100011",
            2447 => "000101000100011",
            2448 => "000101000100011",
            2449 => "000101000100011",
            2450 => "000101000100011",
            2451 => "000101010100100",
            2452 => "000101010100100",
            2453 => "000101010100100",
            2454 => "000101010100100",
            2455 => "000101010100100",
            2456 => "000101010100100",
            2457 => "000101010100100",
            2458 => "000101100101010",
            2459 => "000101100101010",
            2460 => "000101100101010",
            2461 => "000101100101010",
            2462 => "000101100101010",
            2463 => "000101100101010",
            2464 => "000101100101010",
            2465 => "000101110101101",
            2466 => "000101110101101",
            2467 => "000101110101101",
            2468 => "000101110101101",
            2469 => "000101110101101",
            2470 => "000101110101101",
            2471 => "000101110101101",
            2472 => "000110000100010",
            2473 => "000110000100010",
            2474 => "000110000100010",
            2475 => "000110000100010",
            2476 => "000110000100010",
            2477 => "000110000100010",
            2478 => "000110000100010",
            2479 => "000110010100101",
            2480 => "000110010100101",
            2481 => "000110010100101",
            2482 => "000110010100101",
            2483 => "000110010100101",
            2484 => "000110010100101",
            2485 => "000110010100101",
            2486 => "000110100101011",
            2487 => "000110100101011",
            2488 => "000110100101011",
            2489 => "000110100101011",
            2490 => "000110100101011",
            2491 => "000110100101011",
            2492 => "000110100101011",
            2493 => "000110110101100",
            2494 => "000110110101100",
            2495 => "000110110101100",
            2496 => "000110110101100",
            2497 => "000110110101100",
            2498 => "000110110101100",
            2499 => "000110110101100",
            2500 => "000111000101000",
            2501 => "000111000101000",
            2502 => "000111000101000",
            2503 => "000111000101000",
            2504 => "000111000101000",
            2505 => "000111000101000",
            2506 => "000111000101000",
            2507 => "000111010101111",
            2508 => "000111010101111",
            2509 => "000111010101111",
            2510 => "000111010101111",
            2511 => "000111010101111",
            2512 => "000111010101111",
            2513 => "000111010101111",
            2514 => "000111100100001",
            2515 => "000111100100001",
            2516 => "000111100100001",
            2517 => "000111100100001",
            2518 => "000111100100001",
            2519 => "000111100100001",
            2520 => "000111100100001",
            2521 => "000111110100110",
            2522 => "000111110100110",
            2523 => "000111110100110",
            2524 => "000111110100110",
            2525 => "000111110100110",
            2526 => "000111110100110",
            2527 => "000111110100110",
            2528 => "001000000101000",
            2529 => "001000000101000",
            2530 => "001000000101000",
            2531 => "001000000101000",
            2532 => "001000000101000",
            2533 => "001000000101000",
            2534 => "001000000101000",
            2535 => "001000010101111",
            2536 => "001000010101111",
            2537 => "001000010101111",
            2538 => "001000010101111",
            2539 => "001000010101111",
            2540 => "001000010101111",
            2541 => "001000010101111",
            2542 => "001000100100001",
            2543 => "001000100100001",
            2544 => "001000100100001",
            2545 => "001000100100001",
            2546 => "001000100100001",
            2547 => "001000100100001",
            2548 => "001000100100001",
            2549 => "001000110100110",
            2550 => "001000110100110",
            2551 => "001000110100110",
            2552 => "001000110100110",
            2553 => "001000110100110",
            2554 => "001000110100110",
            2555 => "001000110100110",
            2556 => "001001000100010",
            2557 => "001001000100010",
            2558 => "001001000100010",
            2559 => "001001000100010",
            2560 => "001001000100010",
            2561 => "001001000100010",
            2562 => "001001000100010",
            2563 => "001001010100101",
            2564 => "001001010100101",
            2565 => "001001010100101",
            2566 => "001001010100101",
            2567 => "001001010100101",
            2568 => "001001010100101",
            2569 => "001001010100101",
            2570 => "001001100101011",
            2571 => "001001100101011",
            2572 => "001001100101011",
            2573 => "001001100101011",
            2574 => "001001100101011",
            2575 => "001001100101011",
            2576 => "001001100101011",
            2577 => "001001110101100",
            2578 => "001001110101100",
            2579 => "001001110101100",
            2580 => "001001110101100",
            2581 => "001001110101100",
            2582 => "001001110101100",
            2583 => "001001110101100",
            2584 => "001010000100011",
            2585 => "001010000100011",
            2586 => "001010000100011",
            2587 => "001010000100011",
            2588 => "001010000100011",
            2589 => "001010000100011",
            2590 => "001010000100011",
            2591 => "001010010100100",
            2592 => "001010010100100",
            2593 => "001010010100100",
            2594 => "001010010100100",
            2595 => "001010010100100",
            2596 => "001010010100100",
            2597 => "001010010100100",
            2598 => "001010100101010",
            2599 => "001010100101010",
            2600 => "001010100101010",
            2601 => "001010100101010",
            2602 => "001010100101010",
            2603 => "001010100101010",
            2604 => "001010100101010",
            2605 => "001010110101101",
            2606 => "001010110101101",
            2607 => "001010110101101",
            2608 => "001010110101101",
            2609 => "001010110101101",
            2610 => "001010110101101",
            2611 => "001010110101101",
            2612 => "001011000101001",
            2613 => "001011000101001",
            2614 => "001011000101001",
            2615 => "001011000101001",
            2616 => "001011000101001",
            2617 => "001011000101001",
            2618 => "001011000101001",
            2619 => "001011010101110",
            2620 => "001011010101110",
            2621 => "001011010101110",
            2622 => "001011010101110",
            2623 => "001011010101110",
            2624 => "001011010101110",
            2625 => "001011010101110",
            2626 => "001011100100000",
            2627 => "001011100100000",
            2628 => "001011100100000",
            2629 => "001011100100000",
            2630 => "001011100100000",
            2631 => "001011100100000",
            2632 => "001011100100000",
            2633 => "001011110100111",
            2634 => "001011110100111",
            2635 => "001011110100111",
            2636 => "001011110100111",
            2637 => "001011110100111",
            2638 => "001011110100111",
            2639 => "001011110100111",
            2640 => "001100000100100",
            2641 => "001100000100100",
            2642 => "001100000100100",
            2643 => "001100000100100",
            2644 => "001100000100100",
            2645 => "001100000100100",
            2646 => "001100000100100",
            2647 => "001100010100011",
            2648 => "001100010100011",
            2649 => "001100010100011",
            2650 => "001100010100011",
            2651 => "001100010100011",
            2652 => "001100010100011",
            2653 => "001100010100011",
            2654 => "001100100101101",
            2655 => "001100100101101",
            2656 => "001100100101101",
            2657 => "001100100101101",
            2658 => "001100100101101",
            2659 => "001100100101101",
            2660 => "001100100101101",
            2661 => "001100110101010",
            2662 => "001100110101010",
            2663 => "001100110101010",
            2664 => "001100110101010",
            2665 => "001100110101010",
            2666 => "001100110101010",
            2667 => "001100110101010",
            2668 => "001101000101110",
            2669 => "001101000101110",
            2670 => "001101000101110",
            2671 => "001101000101110",
            2672 => "001101000101110",
            2673 => "001101000101110",
            2674 => "001101000101110",
            2675 => "001101010101001",
            2676 => "001101010101001",
            2677 => "001101010101001",
            2678 => "001101010101001",
            2679 => "001101010101001",
            2680 => "001101010101001",
            2681 => "001101010101001",
            2682 => "001101100100111",
            2683 => "001101100100111",
            2684 => "001101100100111",
            2685 => "001101100100111",
            2686 => "001101100100111",
            2687 => "001101100100111",
            2688 => "001101100100111",
            2689 => "001101110100000",
            2690 => "001101110100000",
            2691 => "001101110100000",
            2692 => "001101110100000",
            2693 => "001101110100000",
            2694 => "001101110100000",
            2695 => "001101110100000",
            2696 => "001110000101111",
            2697 => "001110000101111",
            2698 => "001110000101111",
            2699 => "001110000101111",
            2700 => "001110000101111",
            2701 => "001110000101111",
            2702 => "001110000101111",
            2703 => "001110010101000",
            2704 => "001110010101000",
            2705 => "001110010101000",
            2706 => "001110010101000",
            2707 => "001110010101000",
            2708 => "001110010101000",
            2709 => "001110010101000",
            2710 => "001110100100110",
            2711 => "001110100100110",
            2712 => "001110100100110",
            2713 => "001110100100110",
            2714 => "001110100100110",
            2715 => "001110100100110",
            2716 => "001110100100110",
            2717 => "001110110100001",
            2718 => "001110110100001",
            2719 => "001110110100001",
            2720 => "001110110100001",
            2721 => "001110110100001",
            2722 => "001110110100001",
            2723 => "001110110100001",
            2724 => "001111000100101",
            2725 => "001111000100101",
            2726 => "001111000100101",
            2727 => "001111000100101",
            2728 => "001111000100101",
            2729 => "001111000100101",
            2730 => "001111000100101",
            2731 => "001111010100010",
            2732 => "001111010100010",
            2733 => "001111010100010",
            2734 => "001111010100010",
            2735 => "001111010100010",
            2736 => "001111010100010",
            2737 => "001111010100010",
            2738 => "001111100101100",
            2739 => "001111100101100",
            2740 => "001111100101100",
            2741 => "001111100101100",
            2742 => "001111100101100",
            2743 => "001111100101100",
            2744 => "001111100101100",
            2745 => "001111110101011",
            2746 => "001111110101011",
            2747 => "001111110101011",
            2748 => "001111110101011",
            2749 => "001111110101011",
            2750 => "001111110101011",
            2751 => "001111110101011",
            2752 => "010000000101011",
            2753 => "010000000101011",
            2754 => "010000000101011",
            2755 => "010000000101011",
            2756 => "010000000101011",
            2757 => "010000000101011",
            2758 => "010000000101011",
            2759 => "010000010101100",
            2760 => "010000010101100",
            2761 => "010000010101100",
            2762 => "010000010101100",
            2763 => "010000010101100",
            2764 => "010000010101100",
            2765 => "010000010101100",
            2766 => "010000100100010",
            2767 => "010000100100010",
            2768 => "010000100100010",
            2769 => "010000100100010",
            2770 => "010000100100010",
            2771 => "010000100100010",
            2772 => "010000100100010",
            2773 => "010000110100101",
            2774 => "010000110100101",
            2775 => "010000110100101",
            2776 => "010000110100101",
            2777 => "010000110100101",
            2778 => "010000110100101",
            2779 => "010000110100101",
            2780 => "010001000100001",
            2781 => "010001000100001",
            2782 => "010001000100001",
            2783 => "010001000100001",
            2784 => "010001000100001",
            2785 => "010001000100001",
            2786 => "010001000100001",
            2787 => "010001010100110",
            2788 => "010001010100110",
            2789 => "010001010100110",
            2790 => "010001010100110",
            2791 => "010001010100110",
            2792 => "010001010100110",
            2793 => "010001010100110",
            2794 => "010001100101000",
            2795 => "010001100101000",
            2796 => "010001100101000",
            2797 => "010001100101000",
            2798 => "010001100101000",
            2799 => "010001100101000",
            2800 => "010001100101000",
            2801 => "010001110101111",
            2802 => "010001110101111",
            2803 => "010001110101111",
            2804 => "010001110101111",
            2805 => "010001110101111",
            2806 => "010001110101111",
            2807 => "010001110101111",
            2808 => "010010000100000",
            2809 => "010010000100000",
            2810 => "010010000100000",
            2811 => "010010000100000",
            2812 => "010010000100000",
            2813 => "010010000100000",
            2814 => "010010000100000",
            2815 => "010010010100111",
            2816 => "010010010100111",
            2817 => "010010010100111",
            2818 => "010010010100111",
            2819 => "010010010100111",
            2820 => "010010010100111",
            2821 => "010010010100111",
            2822 => "010010100101001",
            2823 => "010010100101001",
            2824 => "010010100101001",
            2825 => "010010100101001",
            2826 => "010010100101001",
            2827 => "010010100101001",
            2828 => "010010100101001",
            2829 => "010010110101110",
            2830 => "010010110101110",
            2831 => "010010110101110",
            2832 => "010010110101110",
            2833 => "010010110101110",
            2834 => "010010110101110",
            2835 => "010010110101110",
            2836 => "010011000101010",
            2837 => "010011000101010",
            2838 => "010011000101010",
            2839 => "010011000101010",
            2840 => "010011000101010",
            2841 => "010011000101010",
            2842 => "010011000101010",
            2843 => "010011010101101",
            2844 => "010011010101101",
            2845 => "010011010101101",
            2846 => "010011010101101",
            2847 => "010011010101101",
            2848 => "010011010101101",
            2849 => "010011010101101",
            2850 => "010011100100011",
            2851 => "010011100100011",
            2852 => "010011100100011",
            2853 => "010011100100011",
            2854 => "010011100100011",
            2855 => "010011100100011",
            2856 => "010011100100011",
            2857 => "010011110100100",
            2858 => "010011110100100",
            2859 => "010011110100100",
            2860 => "010011110100100",
            2861 => "010011110100100",
            2862 => "010011110100100",
            2863 => "010011110100100",
            2864 => "010100000100111",
            2865 => "010100000100111",
            2866 => "010100000100111",
            2867 => "010100000100111",
            2868 => "010100000100111",
            2869 => "010100000100111",
            2870 => "010100000100111",
            2871 => "010100010100000",
            2872 => "010100010100000",
            2873 => "010100010100000",
            2874 => "010100010100000",
            2875 => "010100010100000",
            2876 => "010100010100000",
            2877 => "010100010100000",
            2878 => "010100100101110",
            2879 => "010100100101110",
            2880 => "010100100101110",
            2881 => "010100100101110",
            2882 => "010100100101110",
            2883 => "010100100101110",
            2884 => "010100100101110",
            2885 => "010100110101001",
            2886 => "010100110101001",
            2887 => "010100110101001",
            2888 => "010100110101001",
            2889 => "010100110101001",
            2890 => "010100110101001",
            2891 => "010100110101001",
            2892 => "010101000101101",
            2893 => "010101000101101",
            2894 => "010101000101101",
            2895 => "010101000101101",
            2896 => "010101000101101",
            2897 => "010101000101101",
            2898 => "010101000101101",
            2899 => "010101010101010",
            2900 => "010101010101010",
            2901 => "010101010101010",
            2902 => "010101010101010",
            2903 => "010101010101010",
            2904 => "010101010101010",
            2905 => "010101010101010",
            2906 => "010101100100100",
            2907 => "010101100100100",
            2908 => "010101100100100",
            2909 => "010101100100100",
            2910 => "010101100100100",
            2911 => "010101100100100",
            2912 => "010101100100100",
            2913 => "010101110100011",
            2914 => "010101110100011",
            2915 => "010101110100011",
            2916 => "010101110100011",
            2917 => "010101110100011",
            2918 => "010101110100011",
            2919 => "010101110100011",
            2920 => "010110000101100",
            2921 => "010110000101100",
            2922 => "010110000101100",
            2923 => "010110000101100",
            2924 => "010110000101100",
            2925 => "010110000101100",
            2926 => "010110000101100",
            2927 => "010110010101011",
            2928 => "010110010101011",
            2929 => "010110010101011",
            2930 => "010110010101011",
            2931 => "010110010101011",
            2932 => "010110010101011",
            2933 => "010110010101011",
            2934 => "010110100100101",
            2935 => "010110100100101",
            2936 => "010110100100101",
            2937 => "010110100100101",
            2938 => "010110100100101",
            2939 => "010110100100101",
            2940 => "010110100100101",
            2941 => "010110110100010",
            2942 => "010110110100010",
            2943 => "010110110100010",
            2944 => "010110110100010",
            2945 => "010110110100010",
            2946 => "010110110100010",
            2947 => "010110110100010",
            2948 => "010111000100110",
            2949 => "010111000100110",
            2950 => "010111000100110",
            2951 => "010111000100110",
            2952 => "010111000100110",
            2953 => "010111000100110",
            2954 => "010111000100110",
            2955 => "010111010100001",
            2956 => "010111010100001",
            2957 => "010111010100001",
            2958 => "010111010100001",
            2959 => "010111010100001",
            2960 => "010111010100001",
            2961 => "010111010100001",
            2962 => "010111100101111",
            2963 => "010111100101111",
            2964 => "010111100101111",
            2965 => "010111100101111",
            2966 => "010111100101111",
            2967 => "010111100101111",
            2968 => "010111100101111",
            2969 => "010111110101000",
            2970 => "010111110101000",
            2971 => "010111110101000",
            2972 => "010111110101000",
            2973 => "010111110101000",
            2974 => "010111110101000",
            2975 => "010111110101000",
            2976 => "011000000100110",
            2977 => "011000000100110",
            2978 => "011000000100110",
            2979 => "011000000100110",
            2980 => "011000000100110",
            2981 => "011000000100110",
            2982 => "011000000100110",
            2983 => "011000010100001",
            2984 => "011000010100001",
            2985 => "011000010100001",
            2986 => "011000010100001",
            2987 => "011000010100001",
            2988 => "011000010100001",
            2989 => "011000010100001",
            2990 => "011000100101111",
            2991 => "011000100101111",
            2992 => "011000100101111",
            2993 => "011000100101111",
            2994 => "011000100101111",
            2995 => "011000100101111",
            2996 => "011000100101111",
            2997 => "011000110101000",
            2998 => "011000110101000",
            2999 => "011000110101000",
            3000 => "011000110101000",
            3001 => "011000110101000",
            3002 => "011000110101000",
            3003 => "011000110101000",
            3004 => "011001000101100",
            3005 => "011001000101100",
            3006 => "011001000101100",
            3007 => "011001000101100",
            3008 => "011001000101100",
            3009 => "011001000101100",
            3010 => "011001000101100",
            3011 => "011001010101011",
            3012 => "011001010101011",
            3013 => "011001010101011",
            3014 => "011001010101011",
            3015 => "011001010101011",
            3016 => "011001010101011",
            3017 => "011001010101011",
            3018 => "011001100100101",
            3019 => "011001100100101",
            3020 => "011001100100101",
            3021 => "011001100100101",
            3022 => "011001100100101",
            3023 => "011001100100101",
            3024 => "011001100100101",
            3025 => "011001110100010",
            3026 => "011001110100010",
            3027 => "011001110100010",
            3028 => "011001110100010",
            3029 => "011001110100010",
            3030 => "011001110100010",
            3031 => "011001110100010",
            3032 => "011010000101101",
            3033 => "011010000101101",
            3034 => "011010000101101",
            3035 => "011010000101101",
            3036 => "011010000101101",
            3037 => "011010000101101",
            3038 => "011010000101101",
            3039 => "011010010101010",
            3040 => "011010010101010",
            3041 => "011010010101010",
            3042 => "011010010101010",
            3043 => "011010010101010",
            3044 => "011010010101010",
            3045 => "011010010101010",
            3046 => "011010100100100",
            3047 => "011010100100100",
            3048 => "011010100100100",
            3049 => "011010100100100",
            3050 => "011010100100100",
            3051 => "011010100100100",
            3052 => "011010100100100",
            3053 => "011010110100011",
            3054 => "011010110100011",
            3055 => "011010110100011",
            3056 => "011010110100011",
            3057 => "011010110100011",
            3058 => "011010110100011",
            3059 => "011010110100011",
            3060 => "011011000100111",
            3061 => "011011000100111",
            3062 => "011011000100111",
            3063 => "011011000100111",
            3064 => "011011000100111",
            3065 => "011011000100111",
            3066 => "011011000100111",
            3067 => "011011010100000",
            3068 => "011011010100000",
            3069 => "011011010100000",
            3070 => "011011010100000",
            3071 => "011011010100000",
            3072 => "011011010100000",
            3073 => "011011010100000",
            3074 => "011011100101110",
            3075 => "011011100101110",
            3076 => "011011100101110",
            3077 => "011011100101110",
            3078 => "011011100101110",
            3079 => "011011100101110",
            3080 => "011011100101110",
            3081 => "011011110101001",
            3082 => "011011110101001",
            3083 => "011011110101001",
            3084 => "011011110101001",
            3085 => "011011110101001",
            3086 => "011011110101001",
            3087 => "011011110101001",
            3088 => "011100000101010",
            3089 => "011100000101010",
            3090 => "011100000101010",
            3091 => "011100000101010",
            3092 => "011100000101010",
            3093 => "011100000101010",
            3094 => "011100000101010",
            3095 => "011100010101101",
            3096 => "011100010101101",
            3097 => "011100010101101",
            3098 => "011100010101101",
            3099 => "011100010101101",
            3100 => "011100010101101",
            3101 => "011100010101101",
            3102 => "011100100100011",
            3103 => "011100100100011",
            3104 => "011100100100011",
            3105 => "011100100100011",
            3106 => "011100100100011",
            3107 => "011100100100011",
            3108 => "011100100100011",
            3109 => "011100110100100",
            3110 => "011100110100100",
            3111 => "011100110100100",
            3112 => "011100110100100",
            3113 => "011100110100100",
            3114 => "011100110100100",
            3115 => "011100110100100",
            3116 => "011101000100000",
            3117 => "011101000100000",
            3118 => "011101000100000",
            3119 => "011101000100000",
            3120 => "011101000100000",
            3121 => "011101000100000",
            3122 => "011101000100000",
            3123 => "011101010100111",
            3124 => "011101010100111",
            3125 => "011101010100111",
            3126 => "011101010100111",
            3127 => "011101010100111",
            3128 => "011101010100111",
            3129 => "011101010100111",
            3130 => "011101100101001",
            3131 => "011101100101001",
            3132 => "011101100101001",
            3133 => "011101100101001",
            3134 => "011101100101001",
            3135 => "011101100101001",
            3136 => "011101100101001",
            3137 => "011101110101110",
            3138 => "011101110101110",
            3139 => "011101110101110",
            3140 => "011101110101110",
            3141 => "011101110101110",
            3142 => "011101110101110",
            3143 => "011101110101110",
            3144 => "011110000100001",
            3145 => "011110000100001",
            3146 => "011110000100001",
            3147 => "011110000100001",
            3148 => "011110000100001",
            3149 => "011110000100001",
            3150 => "011110000100001",
            3151 => "011110010100110",
            3152 => "011110010100110",
            3153 => "011110010100110",
            3154 => "011110010100110",
            3155 => "011110010100110",
            3156 => "011110010100110",
            3157 => "011110010100110",
            3158 => "011110100101000",
            3159 => "011110100101000",
            3160 => "011110100101000",
            3161 => "011110100101000",
            3162 => "011110100101000",
            3163 => "011110100101000",
            3164 => "011110100101000",
            3165 => "011110110101111",
            3166 => "011110110101111",
            3167 => "011110110101111",
            3168 => "011110110101111",
            3169 => "011110110101111",
            3170 => "011110110101111",
            3171 => "011110110101111",
            3172 => "011111000101011",
            3173 => "011111000101011",
            3174 => "011111000101011",
            3175 => "011111000101011",
            3176 => "011111000101011",
            3177 => "011111000101011",
            3178 => "011111000101011",
            3179 => "011111010101100",
            3180 => "011111010101100",
            3181 => "011111010101100",
            3182 => "011111010101100",
            3183 => "011111010101100",
            3184 => "011111010101100",
            3185 => "011111010101100",
            3186 => "011111100100010",
            3187 => "011111100100010",
            3188 => "011111100100010",
            3189 => "011111100100010",
            3190 => "011111100100010",
            3191 => "011111100100010",
            3192 => "011111100100010",
            3193 => "011111110100101",
            3194 => "011111110100101",
            3195 => "011111110100101",
            3196 => "011111110100101",
            3197 => "011111110100101",
            3198 => "011111110100101",
            3199 => "011111110100101",
            3200 => "100000000101010",
            3201 => "100000000101010",
            3202 => "100000000101010",
            3203 => "100000000101010",
            3204 => "100000000101010",
            3205 => "100000000101010",
            3206 => "100000000101010",
            3207 => "100000010101101",
            3208 => "100000010101101",
            3209 => "100000010101101",
            3210 => "100000010101101",
            3211 => "100000010101101",
            3212 => "100000010101101",
            3213 => "100000010101101",
            3214 => "100000100100011",
            3215 => "100000100100011",
            3216 => "100000100100011",
            3217 => "100000100100011",
            3218 => "100000100100011",
            3219 => "100000100100011",
            3220 => "100000100100011",
            3221 => "100000110100100",
            3222 => "100000110100100",
            3223 => "100000110100100",
            3224 => "100000110100100",
            3225 => "100000110100100",
            3226 => "100000110100100",
            3227 => "100000110100100",
            3228 => "100001000100000",
            3229 => "100001000100000",
            3230 => "100001000100000",
            3231 => "100001000100000",
            3232 => "100001000100000",
            3233 => "100001000100000",
            3234 => "100001000100000",
            3235 => "100001010100111",
            3236 => "100001010100111",
            3237 => "100001010100111",
            3238 => "100001010100111",
            3239 => "100001010100111",
            3240 => "100001010100111",
            3241 => "100001010100111",
            3242 => "100001100101001",
            3243 => "100001100101001",
            3244 => "100001100101001",
            3245 => "100001100101001",
            3246 => "100001100101001",
            3247 => "100001100101001",
            3248 => "100001100101001",
            3249 => "100001110101110",
            3250 => "100001110101110",
            3251 => "100001110101110",
            3252 => "100001110101110",
            3253 => "100001110101110",
            3254 => "100001110101110",
            3255 => "100001110101110",
            3256 => "100010000100001",
            3257 => "100010000100001",
            3258 => "100010000100001",
            3259 => "100010000100001",
            3260 => "100010000100001",
            3261 => "100010000100001",
            3262 => "100010000100001",
            3263 => "100010010100110",
            3264 => "100010010100110",
            3265 => "100010010100110",
            3266 => "100010010100110",
            3267 => "100010010100110",
            3268 => "100010010100110",
            3269 => "100010010100110",
            3270 => "100010100101000",
            3271 => "100010100101000",
            3272 => "100010100101000",
            3273 => "100010100101000",
            3274 => "100010100101000",
            3275 => "100010100101000",
            3276 => "100010100101000",
            3277 => "100010110101111",
            3278 => "100010110101111",
            3279 => "100010110101111",
            3280 => "100010110101111",
            3281 => "100010110101111",
            3282 => "100010110101111",
            3283 => "100010110101111",
            3284 => "100011000101011",
            3285 => "100011000101011",
            3286 => "100011000101011",
            3287 => "100011000101011",
            3288 => "100011000101011",
            3289 => "100011000101011",
            3290 => "100011000101011",
            3291 => "100011010101100",
            3292 => "100011010101100",
            3293 => "100011010101100",
            3294 => "100011010101100",
            3295 => "100011010101100",
            3296 => "100011010101100",
            3297 => "100011010101100",
            3298 => "100011100100010",
            3299 => "100011100100010",
            3300 => "100011100100010",
            3301 => "100011100100010",
            3302 => "100011100100010",
            3303 => "100011100100010",
            3304 => "100011100100010",
            3305 => "100011110100101",
            3306 => "100011110100101",
            3307 => "100011110100101",
            3308 => "100011110100101",
            3309 => "100011110100101",
            3310 => "100011110100101",
            3311 => "100011110100101",
            3312 => "100100000100110",
            3313 => "100100000100110",
            3314 => "100100000100110",
            3315 => "100100000100110",
            3316 => "100100000100110",
            3317 => "100100000100110",
            3318 => "100100000100110",
            3319 => "100100010100001",
            3320 => "100100010100001",
            3321 => "100100010100001",
            3322 => "100100010100001",
            3323 => "100100010100001",
            3324 => "100100010100001",
            3325 => "100100010100001",
            3326 => "100100100101111",
            3327 => "100100100101111",
            3328 => "100100100101111",
            3329 => "100100100101111",
            3330 => "100100100101111",
            3331 => "100100100101111",
            3332 => "100100100101111",
            3333 => "100100110101000",
            3334 => "100100110101000",
            3335 => "100100110101000",
            3336 => "100100110101000",
            3337 => "100100110101000",
            3338 => "100100110101000",
            3339 => "100100110101000",
            3340 => "100101000101100",
            3341 => "100101000101100",
            3342 => "100101000101100",
            3343 => "100101000101100",
            3344 => "100101000101100",
            3345 => "100101000101100",
            3346 => "100101000101100",
            3347 => "100101010101011",
            3348 => "100101010101011",
            3349 => "100101010101011",
            3350 => "100101010101011",
            3351 => "100101010101011",
            3352 => "100101010101011",
            3353 => "100101010101011",
            3354 => "100101100100101",
            3355 => "100101100100101",
            3356 => "100101100100101",
            3357 => "100101100100101",
            3358 => "100101100100101",
            3359 => "100101100100101",
            3360 => "100101100100101",
            3361 => "100101110100010",
            3362 => "100101110100010",
            3363 => "100101110100010",
            3364 => "100101110100010",
            3365 => "100101110100010",
            3366 => "100101110100010",
            3367 => "100101110100010",
            3368 => "100110000101101",
            3369 => "100110000101101",
            3370 => "100110000101101",
            3371 => "100110000101101",
            3372 => "100110000101101",
            3373 => "100110000101101",
            3374 => "100110000101101",
            3375 => "100110010101010",
            3376 => "100110010101010",
            3377 => "100110010101010",
            3378 => "100110010101010",
            3379 => "100110010101010",
            3380 => "100110010101010",
            3381 => "100110010101010",
            3382 => "100110100100100",
            3383 => "100110100100100",
            3384 => "100110100100100",
            3385 => "100110100100100",
            3386 => "100110100100100",
            3387 => "100110100100100",
            3388 => "100110100100100",
            3389 => "100110110100011",
            3390 => "100110110100011",
            3391 => "100110110100011",
            3392 => "100110110100011",
            3393 => "100110110100011",
            3394 => "100110110100011",
            3395 => "100110110100011",
            3396 => "100111000100111",
            3397 => "100111000100111",
            3398 => "100111000100111",
            3399 => "100111000100111",
            3400 => "100111000100111",
            3401 => "100111000100111",
            3402 => "100111000100111",
            3403 => "100111010100000",
            3404 => "100111010100000",
            3405 => "100111010100000",
            3406 => "100111010100000",
            3407 => "100111010100000",
            3408 => "100111010100000",
            3409 => "100111010100000",
            3410 => "100111100101110",
            3411 => "100111100101110",
            3412 => "100111100101110",
            3413 => "100111100101110",
            3414 => "100111100101110",
            3415 => "100111100101110",
            3416 => "100111100101110",
            3417 => "100111110101001",
            3418 => "100111110101001",
            3419 => "100111110101001",
            3420 => "100111110101001",
            3421 => "100111110101001",
            3422 => "100111110101001",
            3423 => "100111110101001",
            3424 => "101000000100111",
            3425 => "101000000100111",
            3426 => "101000000100111",
            3427 => "101000000100111",
            3428 => "101000000100111",
            3429 => "101000000100111",
            3430 => "101000000100111",
            3431 => "101000010100000",
            3432 => "101000010100000",
            3433 => "101000010100000",
            3434 => "101000010100000",
            3435 => "101000010100000",
            3436 => "101000010100000",
            3437 => "101000010100000",
            3438 => "101000100101110",
            3439 => "101000100101110",
            3440 => "101000100101110",
            3441 => "101000100101110",
            3442 => "101000100101110",
            3443 => "101000100101110",
            3444 => "101000100101110",
            3445 => "101000110101001",
            3446 => "101000110101001",
            3447 => "101000110101001",
            3448 => "101000110101001",
            3449 => "101000110101001",
            3450 => "101000110101001",
            3451 => "101000110101001",
            3452 => "101001000101101",
            3453 => "101001000101101",
            3454 => "101001000101101",
            3455 => "101001000101101",
            3456 => "101001000101101",
            3457 => "101001000101101",
            3458 => "101001000101101",
            3459 => "101001010101010",
            3460 => "101001010101010",
            3461 => "101001010101010",
            3462 => "101001010101010",
            3463 => "101001010101010",
            3464 => "101001010101010",
            3465 => "101001010101010",
            3466 => "101001100100100",
            3467 => "101001100100100",
            3468 => "101001100100100",
            3469 => "101001100100100",
            3470 => "101001100100100",
            3471 => "101001100100100",
            3472 => "101001100100100",
            3473 => "101001110100011",
            3474 => "101001110100011",
            3475 => "101001110100011",
            3476 => "101001110100011",
            3477 => "101001110100011",
            3478 => "101001110100011",
            3479 => "101001110100011",
            3480 => "101010000101100",
            3481 => "101010000101100",
            3482 => "101010000101100",
            3483 => "101010000101100",
            3484 => "101010000101100",
            3485 => "101010000101100",
            3486 => "101010000101100",
            3487 => "101010010101011",
            3488 => "101010010101011",
            3489 => "101010010101011",
            3490 => "101010010101011",
            3491 => "101010010101011",
            3492 => "101010010101011",
            3493 => "101010010101011",
            3494 => "101010100100101",
            3495 => "101010100100101",
            3496 => "101010100100101",
            3497 => "101010100100101",
            3498 => "101010100100101",
            3499 => "101010100100101",
            3500 => "101010100100101",
            3501 => "101010110100010",
            3502 => "101010110100010",
            3503 => "101010110100010",
            3504 => "101010110100010",
            3505 => "101010110100010",
            3506 => "101010110100010",
            3507 => "101010110100010",
            3508 => "101011000100110",
            3509 => "101011000100110",
            3510 => "101011000100110",
            3511 => "101011000100110",
            3512 => "101011000100110",
            3513 => "101011000100110",
            3514 => "101011000100110",
            3515 => "101011010100001",
            3516 => "101011010100001",
            3517 => "101011010100001",
            3518 => "101011010100001",
            3519 => "101011010100001",
            3520 => "101011010100001",
            3521 => "101011010100001",
            3522 => "101011100101111",
            3523 => "101011100101111",
            3524 => "101011100101111",
            3525 => "101011100101111",
            3526 => "101011100101111",
            3527 => "101011100101111",
            3528 => "101011100101111",
            3529 => "101011110101000",
            3530 => "101011110101000",
            3531 => "101011110101000",
            3532 => "101011110101000",
            3533 => "101011110101000",
            3534 => "101011110101000",
            3535 => "101011110101000",
            3536 => "101100000101011",
            3537 => "101100000101011",
            3538 => "101100000101011",
            3539 => "101100000101011",
            3540 => "101100000101011",
            3541 => "101100000101011",
            3542 => "101100000101011",
            3543 => "101100010101100",
            3544 => "101100010101100",
            3545 => "101100010101100",
            3546 => "101100010101100",
            3547 => "101100010101100",
            3548 => "101100010101100",
            3549 => "101100010101100",
            3550 => "101100100100010",
            3551 => "101100100100010",
            3552 => "101100100100010",
            3553 => "101100100100010",
            3554 => "101100100100010",
            3555 => "101100100100010",
            3556 => "101100100100010",
            3557 => "101100110100101",
            3558 => "101100110100101",
            3559 => "101100110100101",
            3560 => "101100110100101",
            3561 => "101100110100101",
            3562 => "101100110100101",
            3563 => "101100110100101",
            3564 => "101101000100001",
            3565 => "101101000100001",
            3566 => "101101000100001",
            3567 => "101101000100001",
            3568 => "101101000100001",
            3569 => "101101000100001",
            3570 => "101101000100001",
            3571 => "101101010100110",
            3572 => "101101010100110",
            3573 => "101101010100110",
            3574 => "101101010100110",
            3575 => "101101010100110",
            3576 => "101101010100110",
            3577 => "101101010100110",
            3578 => "101101100101000",
            3579 => "101101100101000",
            3580 => "101101100101000",
            3581 => "101101100101000",
            3582 => "101101100101000",
            3583 => "101101100101000",
            3584 => "101101100101000",
            3585 => "101101110101111",
            3586 => "101101110101111",
            3587 => "101101110101111",
            3588 => "101101110101111",
            3589 => "101101110101111",
            3590 => "101101110101111",
            3591 => "101101110101111",
            3592 => "101110000100000",
            3593 => "101110000100000",
            3594 => "101110000100000",
            3595 => "101110000100000",
            3596 => "101110000100000",
            3597 => "101110000100000",
            3598 => "101110000100000",
            3599 => "101110010100111",
            3600 => "101110010100111",
            3601 => "101110010100111",
            3602 => "101110010100111",
            3603 => "101110010100111",
            3604 => "101110010100111",
            3605 => "101110010100111",
            3606 => "101110100101001",
            3607 => "101110100101001",
            3608 => "101110100101001",
            3609 => "101110100101001",
            3610 => "101110100101001",
            3611 => "101110100101001",
            3612 => "101110100101001",
            3613 => "101110110101110",
            3614 => "101110110101110",
            3615 => "101110110101110",
            3616 => "101110110101110",
            3617 => "101110110101110",
            3618 => "101110110101110",
            3619 => "101110110101110",
            3620 => "101111000101010",
            3621 => "101111000101010",
            3622 => "101111000101010",
            3623 => "101111000101010",
            3624 => "101111000101010",
            3625 => "101111000101010",
            3626 => "101111000101010",
            3627 => "101111010101101",
            3628 => "101111010101101",
            3629 => "101111010101101",
            3630 => "101111010101101",
            3631 => "101111010101101",
            3632 => "101111010101101",
            3633 => "101111010101101",
            3634 => "101111100100011",
            3635 => "101111100100011",
            3636 => "101111100100011",
            3637 => "101111100100011",
            3638 => "101111100100011",
            3639 => "101111100100011",
            3640 => "101111100100011",
            3641 => "101111110100100",
            3642 => "101111110100100",
            3643 => "101111110100100",
            3644 => "101111110100100",
            3645 => "101111110100100",
            3646 => "101111110100100",
            3647 => "101111110100100",
            3648 => "110000000100100",
            3649 => "110000000100100",
            3650 => "110000000100100",
            3651 => "110000000100100",
            3652 => "110000000100100",
            3653 => "110000000100100",
            3654 => "110000000100100",
            3655 => "110000010100011",
            3656 => "110000010100011",
            3657 => "110000010100011",
            3658 => "110000010100011",
            3659 => "110000010100011",
            3660 => "110000010100011",
            3661 => "110000010100011",
            3662 => "110000100101101",
            3663 => "110000100101101",
            3664 => "110000100101101",
            3665 => "110000100101101",
            3666 => "110000100101101",
            3667 => "110000100101101",
            3668 => "110000100101101",
            3669 => "110000110101010",
            3670 => "110000110101010",
            3671 => "110000110101010",
            3672 => "110000110101010",
            3673 => "110000110101010",
            3674 => "110000110101010",
            3675 => "110000110101010",
            3676 => "110001000101110",
            3677 => "110001000101110",
            3678 => "110001000101110",
            3679 => "110001000101110",
            3680 => "110001000101110",
            3681 => "110001000101110",
            3682 => "110001000101110",
            3683 => "110001010101001",
            3684 => "110001010101001",
            3685 => "110001010101001",
            3686 => "110001010101001",
            3687 => "110001010101001",
            3688 => "110001010101001",
            3689 => "110001010101001",
            3690 => "110001100100111",
            3691 => "110001100100111",
            3692 => "110001100100111",
            3693 => "110001100100111",
            3694 => "110001100100111",
            3695 => "110001100100111",
            3696 => "110001100100111",
            3697 => "110001110100000",
            3698 => "110001110100000",
            3699 => "110001110100000",
            3700 => "110001110100000",
            3701 => "110001110100000",
            3702 => "110001110100000",
            3703 => "110001110100000",
            3704 => "110010000101111",
            3705 => "110010000101111",
            3706 => "110010000101111",
            3707 => "110010000101111",
            3708 => "110010000101111",
            3709 => "110010000101111",
            3710 => "110010000101111",
            3711 => "110010010101000",
            3712 => "110010010101000",
            3713 => "110010010101000",
            3714 => "110010010101000",
            3715 => "110010010101000",
            3716 => "110010010101000",
            3717 => "110010010101000",
            3718 => "110010100100110",
            3719 => "110010100100110",
            3720 => "110010100100110",
            3721 => "110010100100110",
            3722 => "110010100100110",
            3723 => "110010100100110",
            3724 => "110010100100110",
            3725 => "110010110100001",
            3726 => "110010110100001",
            3727 => "110010110100001",
            3728 => "110010110100001",
            3729 => "110010110100001",
            3730 => "110010110100001",
            3731 => "110010110100001",
            3732 => "110011000100101",
            3733 => "110011000100101",
            3734 => "110011000100101",
            3735 => "110011000100101",
            3736 => "110011000100101",
            3737 => "110011000100101",
            3738 => "110011000100101",
            3739 => "110011010100010",
            3740 => "110011010100010",
            3741 => "110011010100010",
            3742 => "110011010100010",
            3743 => "110011010100010",
            3744 => "110011010100010",
            3745 => "110011010100010",
            3746 => "110011100101100",
            3747 => "110011100101100",
            3748 => "110011100101100",
            3749 => "110011100101100",
            3750 => "110011100101100",
            3751 => "110011100101100",
            3752 => "110011100101100",
            3753 => "110011110101011",
            3754 => "110011110101011",
            3755 => "110011110101011",
            3756 => "110011110101011",
            3757 => "110011110101011",
            3758 => "110011110101011",
            3759 => "110011110101011",
            3760 => "110100000101000",
            3761 => "110100000101000",
            3762 => "110100000101000",
            3763 => "110100000101000",
            3764 => "110100000101000",
            3765 => "110100000101000",
            3766 => "110100000101000",
            3767 => "110100010101111",
            3768 => "110100010101111",
            3769 => "110100010101111",
            3770 => "110100010101111",
            3771 => "110100010101111",
            3772 => "110100010101111",
            3773 => "110100010101111",
            3774 => "110100100100001",
            3775 => "110100100100001",
            3776 => "110100100100001",
            3777 => "110100100100001",
            3778 => "110100100100001",
            3779 => "110100100100001",
            3780 => "110100100100001",
            3781 => "110100110100110",
            3782 => "110100110100110",
            3783 => "110100110100110",
            3784 => "110100110100110",
            3785 => "110100110100110",
            3786 => "110100110100110",
            3787 => "110100110100110",
            3788 => "110101000100010",
            3789 => "110101000100010",
            3790 => "110101000100010",
            3791 => "110101000100010",
            3792 => "110101000100010",
            3793 => "110101000100010",
            3794 => "110101000100010",
            3795 => "110101010100101",
            3796 => "110101010100101",
            3797 => "110101010100101",
            3798 => "110101010100101",
            3799 => "110101010100101",
            3800 => "110101010100101",
            3801 => "110101010100101",
            3802 => "110101100101011",
            3803 => "110101100101011",
            3804 => "110101100101011",
            3805 => "110101100101011",
            3806 => "110101100101011",
            3807 => "110101100101011",
            3808 => "110101100101011",
            3809 => "110101110101100",
            3810 => "110101110101100",
            3811 => "110101110101100",
            3812 => "110101110101100",
            3813 => "110101110101100",
            3814 => "110101110101100",
            3815 => "110101110101100",
            3816 => "110110000100011",
            3817 => "110110000100011",
            3818 => "110110000100011",
            3819 => "110110000100011",
            3820 => "110110000100011",
            3821 => "110110000100011",
            3822 => "110110000100011",
            3823 => "110110010100100",
            3824 => "110110010100100",
            3825 => "110110010100100",
            3826 => "110110010100100",
            3827 => "110110010100100",
            3828 => "110110010100100",
            3829 => "110110010100100",
            3830 => "110110100101010",
            3831 => "110110100101010",
            3832 => "110110100101010",
            3833 => "110110100101010",
            3834 => "110110100101010",
            3835 => "110110100101010",
            3836 => "110110100101010",
            3837 => "110110110101101",
            3838 => "110110110101101",
            3839 => "110110110101101",
            3840 => "110110110101101",
            3841 => "110110110101101",
            3842 => "110110110101101",
            3843 => "110110110101101",
            3844 => "110111000101001",
            3845 => "110111000101001",
            3846 => "110111000101001",
            3847 => "110111000101001",
            3848 => "110111000101001",
            3849 => "110111000101001",
            3850 => "110111000101001",
            3851 => "110111010101110",
            3852 => "110111010101110",
            3853 => "110111010101110",
            3854 => "110111010101110",
            3855 => "110111010101110",
            3856 => "110111010101110",
            3857 => "110111010101110",
            3858 => "110111100100000",
            3859 => "110111100100000",
            3860 => "110111100100000",
            3861 => "110111100100000",
            3862 => "110111100100000",
            3863 => "110111100100000",
            3864 => "110111100100000",
            3865 => "110111110100111",
            3866 => "110111110100111",
            3867 => "110111110100111",
            3868 => "110111110100111",
            3869 => "110111110100111",
            3870 => "110111110100111",
            3871 => "110111110100111",
            3872 => "111000000101001",
            3873 => "111000000101001",
            3874 => "111000000101001",
            3875 => "111000000101001",
            3876 => "111000000101001",
            3877 => "111000000101001",
            3878 => "111000000101001",
            3879 => "111000010101110",
            3880 => "111000010101110",
            3881 => "111000010101110",
            3882 => "111000010101110",
            3883 => "111000010101110",
            3884 => "111000010101110",
            3885 => "111000010101110",
            3886 => "111000100100000",
            3887 => "111000100100000",
            3888 => "111000100100000",
            3889 => "111000100100000",
            3890 => "111000100100000",
            3891 => "111000100100000",
            3892 => "111000100100000",
            3893 => "111000110100111",
            3894 => "111000110100111",
            3895 => "111000110100111",
            3896 => "111000110100111",
            3897 => "111000110100111",
            3898 => "111000110100111",
            3899 => "111000110100111",
            3900 => "111001000100011",
            3901 => "111001000100011",
            3902 => "111001000100011",
            3903 => "111001000100011",
            3904 => "111001000100011",
            3905 => "111001000100011",
            3906 => "111001000100011",
            3907 => "111001010100100",
            3908 => "111001010100100",
            3909 => "111001010100100",
            3910 => "111001010100100",
            3911 => "111001010100100",
            3912 => "111001010100100",
            3913 => "111001010100100",
            3914 => "111001100101010",
            3915 => "111001100101010",
            3916 => "111001100101010",
            3917 => "111001100101010",
            3918 => "111001100101010",
            3919 => "111001100101010",
            3920 => "111001100101010",
            3921 => "111001110101101",
            3922 => "111001110101101",
            3923 => "111001110101101",
            3924 => "111001110101101",
            3925 => "111001110101101",
            3926 => "111001110101101",
            3927 => "111001110101101",
            3928 => "111010000100010",
            3929 => "111010000100010",
            3930 => "111010000100010",
            3931 => "111010000100010",
            3932 => "111010000100010",
            3933 => "111010000100010",
            3934 => "111010000100010",
            3935 => "111010010100101",
            3936 => "111010010100101",
            3937 => "111010010100101",
            3938 => "111010010100101",
            3939 => "111010010100101",
            3940 => "111010010100101",
            3941 => "111010010100101",
            3942 => "111010100101011",
            3943 => "111010100101011",
            3944 => "111010100101011",
            3945 => "111010100101011",
            3946 => "111010100101011",
            3947 => "111010100101011",
            3948 => "111010100101011",
            3949 => "111010110101100",
            3950 => "111010110101100",
            3951 => "111010110101100",
            3952 => "111010110101100",
            3953 => "111010110101100",
            3954 => "111010110101100",
            3955 => "111010110101100",
            3956 => "111011000101000",
            3957 => "111011000101000",
            3958 => "111011000101000",
            3959 => "111011000101000",
            3960 => "111011000101000",
            3961 => "111011000101000",
            3962 => "111011000101000",
            3963 => "111011010101111",
            3964 => "111011010101111",
            3965 => "111011010101111",
            3966 => "111011010101111",
            3967 => "111011010101111",
            3968 => "111011010101111",
            3969 => "111011010101111",
            3970 => "111011100100001",
            3971 => "111011100100001",
            3972 => "111011100100001",
            3973 => "111011100100001",
            3974 => "111011100100001",
            3975 => "111011100100001",
            3976 => "111011100100001",
            3977 => "111011110100110",
            3978 => "111011110100110",
            3979 => "111011110100110",
            3980 => "111011110100110",
            3981 => "111011110100110",
            3982 => "111011110100110",
            3983 => "111011110100110",
            3984 => "111100000100101",
            3985 => "111100000100101",
            3986 => "111100000100101",
            3987 => "111100000100101",
            3988 => "111100000100101",
            3989 => "111100000100101",
            3990 => "111100000100101",
            3991 => "111100010100010",
            3992 => "111100010100010",
            3993 => "111100010100010",
            3994 => "111100010100010",
            3995 => "111100010100010",
            3996 => "111100010100010",
            3997 => "111100010100010",
            3998 => "111100100101100",
            3999 => "111100100101100",
            4000 => "111100100101100",
            4001 => "111100100101100",
            4002 => "111100100101100",
            4003 => "111100100101100",
            4004 => "111100100101100",
            4005 => "111100110101011",
            4006 => "111100110101011",
            4007 => "111100110101011",
            4008 => "111100110101011",
            4009 => "111100110101011",
            4010 => "111100110101011",
            4011 => "111100110101011",
            4012 => "111101000101111",
            4013 => "111101000101111",
            4014 => "111101000101111",
            4015 => "111101000101111",
            4016 => "111101000101111",
            4017 => "111101000101111",
            4018 => "111101000101111",
            4019 => "111101010101000",
            4020 => "111101010101000",
            4021 => "111101010101000",
            4022 => "111101010101000",
            4023 => "111101010101000",
            4024 => "111101010101000",
            4025 => "111101010101000",
            4026 => "111101100100110",
            4027 => "111101100100110",
            4028 => "111101100100110",
            4029 => "111101100100110",
            4030 => "111101100100110",
            4031 => "111101100100110",
            4032 => "111101100100110",
            4033 => "111101110100001",
            4034 => "111101110100001",
            4035 => "111101110100001",
            4036 => "111101110100001",
            4037 => "111101110100001",
            4038 => "111101110100001",
            4039 => "111101110100001",
            4040 => "111110000101110",
            4041 => "111110000101110",
            4042 => "111110000101110",
            4043 => "111110000101110",
            4044 => "111110000101110",
            4045 => "111110000101110",
            4046 => "111110000101110",
            4047 => "111110010101001",
            4048 => "111110010101001",
            4049 => "111110010101001",
            4050 => "111110010101001",
            4051 => "111110010101001",
            4052 => "111110010101001",
            4053 => "111110010101001",
            4054 => "111110100100111",
            4055 => "111110100100111",
            4056 => "111110100100111",
            4057 => "111110100100111",
            4058 => "111110100100111",
            4059 => "111110100100111",
            4060 => "111110100100111",
            4061 => "111110110100000",
            4062 => "111110110100000",
            4063 => "111110110100000",
            4064 => "111110110100000",
            4065 => "111110110100000",
            4066 => "111110110100000",
            4067 => "111110110100000",
            4068 => "111111000100100",
            4069 => "111111000100100",
            4070 => "111111000100100",
            4071 => "111111000100100",
            4072 => "111111000100100",
            4073 => "111111000100100",
            4074 => "111111000100100",
            4075 => "111111010100011",
            4076 => "111111010100011",
            4077 => "111111010100011",
            4078 => "111111010100011",
            4079 => "111111010100011",
            4080 => "111111010100011",
            4081 => "111111010100011",
            4082 => "111111100101101",
            4083 => "111111100101101",
            4084 => "111111100101101",
            4085 => "111111100101101",
            4086 => "111111100101101",
            4087 => "111111100101101",
            4088 => "111111100101101",
            4089 => "111111110101010",
            4090 => "111111110101010",
            4091 => "111111110101010",
            4092 => "111111110101010",
            4093 => "111111110101010",
            4094 => "111111110101010",
            4095 => "111111110101010"
	);
end package;
