library ieee;
use ieee.std_logic_1164.all;

use work.liaison_tb_data.all;
use work.txt_util.all;

entity liaison_tb is
end liaison_tb;

architecture tb_arch of liaison_tb is
	-- Component declaration of the tested unit
	component liaison
	port(
		clk : in STD_LOGIC;
		mp_data : in STD_LOGIC_VECTOR(3 downto 0);
		reset : in STD_LOGIC;
		di_ready : in STD_LOGIC;
		do_ready : out STD_LOGIC;
		voted_data : out STD_LOGIC );
	end component;
	
	signal clk_period : time := 40 ns;
	
	-- Stimulus signals - signals mapped to the input and inout ports of tested entity
	signal clk : STD_LOGIC;
	signal mp_data : STD_LOGIC_VECTOR(3 downto 0);
	signal reset : STD_LOGIC;
	signal di_ready : STD_LOGIC;   
	
	-- Observed signals - signals mapped to the output ports of tested entity
	signal do_ready : STD_LOGIC;
	signal voted_data : STD_LOGIC;

begin
	process begin
	    clk <= '1';
	    wait for clk_period/2;
	    clk <= '0';
	    wait for clk_period/2;
	end process;
	
	-- Unit Under Test port map
	UUT : liaison
		port map (
			clk => clk,
			mp_data => mp_data,
			reset => reset,
			di_ready => di_ready,
			do_ready => do_ready,
			voted_data => voted_data
		);
 
	
	-- Feed autogenerated test vectors into the system
	-- The vectors have the following strucutre:
	-- 0 => (
	--      0 => "10111010", -- MCU 0 input
	--	    1 => "10111010", -- MCU 1 input
	--	    2 => "10111010", -- MCU 2 input
	--	    3 => "10111010", -- MCU 3 input
	--      4 => "--------"  -- Reset, either 1's or 0's -> 1's the system is reset 
	--                                 before this input
	-- ),
	
	input_process: process begin
	    assert false report "Liaison TB: input start" severity note;
	    	    
		for i in input'range loop
		
		    if input(i, 4)(0) = '1' then		        
		        assert false report "Resetting before input #"&str(i);
		        
		        -- Wait for 8 periods, to make sure any output has completed, then reset
		        if i /= 0 then wait for clk_period*8; end if;
	            reset <= '1';
	            wait for clk_period*2;
	            wait until falling_edge(clk);
	            reset <= '0';
	        end if;
		    		    
		    for j in input(i, 0)'range loop		        
		        if j = 7 then	            
        		    di_ready <= '1';
        		else 
        		    di_ready <= '0';
        		end if;
		        -- Input is an array of test cases, each test is an array of four inputs, and
		        -- each input is a vector of bits. input(i, j, k) test i, MCU j, bit # k.
		        mp_data <= input(i, 0)(j) & input(i, 1)(j) & input(i, 2)(j) & input(i, 3)(j);
		        
		        wait until falling_edge(clk);
		    end loop;
		    
		    -- min 15 cycle between inputs, 15-7 = 8
		    wait for clk_period*8;
		    wait until falling_edge(clk);
		    assert false report "Input #"&str(i)&" done";
		end loop;
		
		assert false report "Liaison TB: input complete" severity note;
		wait;
	end process;
	
	-- Output verification process
	-- Tests the output of the system against a array of autogenerated output vectors
	verification_process: process 
	    variable actual_output : std_logic_vector(14 downto 0) := "000000000000000";
	    variable errors : integer := 0;
	begin
	    for i in output'range loop
		    -- wait for output signal signal to be toggled
		    wait until rising_edge(do_ready);
		    -- Then for the falling edge, as this is when the external system samples
		    wait until falling_edge(clk);
		    
		    -- Build a actual output vector
		    for j in output(i)'range loop
		        actual_output(j) := voted_data;	
		        wait until falling_edge(clk);
		    end loop;
		    		    
		    -- Compare actual and expected output
		    if actual_output = output(i) then
		        assert false report "Output "&str(i)&": OK";
		    else 
    		    assert false report "Output "&str(i)&": Expected " & str(output(i)) & " got " & str(actual_output) severity error;
    		    errors := errors + 1;
    		end if;
		end loop;
		
		if errors = 0 then
		    report "VERIFICATION SUCCESSFULL" severity note;
		else 
            report "VERIFICATION FAILED WITH "&str(errors)&" error(s)" severity failure;
        end if;
        
		wait;
	end process;
end tb_arch;
